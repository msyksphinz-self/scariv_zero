package riscv_vec_conf_pkg;

  parameter VLEN_W = 256;
  parameter DLEN_W = 256;

endpackage // riscv_vec_pkg
