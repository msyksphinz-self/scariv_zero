package recurse_pkg;

localparam MAX = 0;

endpackage // recurse_pkg
