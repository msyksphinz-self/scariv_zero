package riscv_fpu_pkg;

parameter FLEN_W = 64;

endpackage // riscv_fpu_pkg
