package msrh_ic_pkg;

typedef enum logic [ 1: 0] {
  ICInit,
  ICReq,
  ICInvalidate,
  ICResp
} ic_state_t;


endpackage // msrh_ic_pkg
