package riscv_vec_conf_pkg;

  parameter VLEN_W = 0;
  parameter DLEN_W = 0;

endpackage // riscv_vec_pkg
