module msrh_bru_pipe
  import decoder_bru_ctrl_pkg::*;
#(
  parameter RV_ENTRY_SIZE = 32
  )
(
  input logic                       i_clk,
  input logic                       i_reset_n,

  input                             msrh_pkg::issue_t rv0_issue,
  input logic [RV_ENTRY_SIZE-1:0]   rv0_index,
  input                             msrh_pkg::phy_wr_t ex1_i_phy_wr[msrh_pkg::TGT_BUS_SIZE],

  // Commit notification
  input msrh_pkg::commit_blk_t      i_commit,

  input msrh_pkg::mispred_t         i_mispred_lsu[msrh_conf_pkg::LSU_INST_NUM],

 regread_if.master ex1_regread_rs1,
 regread_if.master ex1_regread_rs2,

  output                            msrh_pkg::early_wr_t o_ex1_early_wr,
  output                            msrh_pkg::phy_wr_t o_ex3_phy_wr,

  done_if.master   ex3_done_if,
  br_upd_if.master ex3_br_upd_if
);

typedef struct packed {
  op_t  op;
  imm_t imm;
  logic wr_rd;
} pipe_ctrl_t;

logic   w_commit_flushed;

msrh_pkg::issue_t                        r_ex0_issue;
logic [RV_ENTRY_SIZE-1: 0] w_ex0_index;
pipe_ctrl_t                              w_ex0_pipe_ctrl;
logic                      w_ex0_br_flush;

pipe_ctrl_t                              r_ex1_pipe_ctrl;
msrh_pkg::issue_t                        r_ex1_issue;
msrh_pkg::issue_t                        w_ex1_issue_next;
logic [RV_ENTRY_SIZE-1: 0] r_ex1_index;
logic                      w_ex1_br_flush;
logic                      r_ex1_dead;

logic [msrh_pkg::TGT_BUS_SIZE-1:0] w_ex2_rs1_fwd_valid;
logic [msrh_pkg::TGT_BUS_SIZE-1:0] w_ex2_rs2_fwd_valid;
riscv_pkg::xlen_t w_ex2_tgt_data          [msrh_pkg::TGT_BUS_SIZE];
riscv_pkg::xlen_t w_ex2_rs1_fwd_data;
riscv_pkg::xlen_t w_ex2_rs2_fwd_data;

riscv_pkg::xlen_t w_ex2_rs1_selected_data;
riscv_pkg::xlen_t w_ex2_rs2_selected_data;

logic                                    w_ex2_rs1_pred_hit;
logic                                    w_ex2_rs2_pred_hit;

logic                                    w_ex1_rs1_lsu_mispred;
logic                                    w_ex1_rs2_lsu_mispred;
logic                                    w_ex1_rs1_mispred;
logic                                    w_ex1_rs2_mispred;

pipe_ctrl_t                              r_ex2_pipe_ctrl;
msrh_pkg::issue_t                        r_ex2_issue;
msrh_pkg::issue_t                        w_ex2_issue_next;
logic [RV_ENTRY_SIZE-1: 0]               r_ex2_index;
riscv_pkg::xlen_t            r_ex2_rs1_data;
riscv_pkg::xlen_t            r_ex2_rs2_data;
logic [riscv_pkg::VADDR_W-1: 0]          w_ex2_br_vaddr;
logic                                    r_ex2_wr_valid;
logic                                    w_ex2_br_flush;
logic                                    r_ex2_dead;

msrh_pkg::issue_t                        r_ex3_issue;
msrh_pkg::issue_t                        w_ex3_issue_next;
pipe_ctrl_t                              r_ex3_pipe_ctrl;
logic                                    r_ex3_result;
logic [RV_ENTRY_SIZE-1: 0]               r_ex3_index;
logic [riscv_pkg::VADDR_W-1: 0]          r_ex3_br_vaddr;
logic                                    r_ex3_rs1_pred_hit;
logic                                    r_ex3_rs2_pred_hit;
logic                                    r_ex3_dead;

always_comb begin
  r_ex0_issue = rv0_issue;
  w_ex0_index = rv0_index;
end

decoder_bru_ctrl u_pipe_ctrl (
  .inst(r_ex0_issue.inst),
  .op  (w_ex0_pipe_ctrl.op),
  .imm (w_ex0_pipe_ctrl.imm),
  .wr_rd (w_ex0_pipe_ctrl.wr_rd)
);

assign ex1_regread_rs1.valid = r_ex1_issue.valid & r_ex1_issue.rd_regs[0].valid;
assign ex1_regread_rs1.rnid  = r_ex1_issue.rd_regs[0].rnid;

assign ex1_regread_rs2.valid = r_ex1_issue.valid & r_ex1_issue.rd_regs[1].valid;
assign ex1_regread_rs2.rnid  = r_ex1_issue.rd_regs[1].rnid;

// EX0 brtag flush check
assign w_ex0_br_flush  = msrh_pkg::is_br_flush_target(r_ex0_issue.br_mask, ex3_br_upd_if.brtag,
                                                      ex3_br_upd_if.dead, ex3_br_upd_if.mispredict) & ex3_br_upd_if.update & r_ex0_issue.valid;

always_comb begin
  w_ex1_issue_next = r_ex0_issue;
end

always_ff @(posedge i_clk, negedge i_reset_n) begin
  if (!i_reset_n) begin
    r_ex1_issue <= 'h0;
    r_ex1_index <= 'h0;
    r_ex1_pipe_ctrl <= 'h0;
    r_ex1_dead <= 1'b0;
  end else begin
    r_ex1_issue <= r_ex0_issue;
    r_ex1_index <= w_ex0_index;
    r_ex1_pipe_ctrl <= w_ex0_pipe_ctrl;
    r_ex1_dead <= r_ex0_issue.valid & (w_ex0_br_flush | w_commit_flushed);
  end
end

select_mispred_bus rs1_mispred_select
(
 .i_entry_rnid (r_ex1_issue.rd_regs[0].rnid),
 .i_entry_type (r_ex1_issue.rd_regs[0].typ),
 .i_mispred    (i_mispred_lsu),

 .o_mispred    (w_ex1_rs1_lsu_mispred)
 );


select_mispred_bus rs2_mispred_select
(
 .i_entry_rnid (r_ex1_issue.rd_regs[1].rnid),
 .i_entry_type (r_ex1_issue.rd_regs[1].typ),
 .i_mispred    (i_mispred_lsu),

 .o_mispred    (w_ex1_rs2_lsu_mispred)
 );

assign w_commit_flushed = msrh_pkg::is_flushed_commit(i_commit);


assign w_ex1_rs1_mispred = r_ex1_issue.rd_regs[0].valid & r_ex1_issue.rd_regs[0].predict_ready ? w_ex1_rs1_lsu_mispred : 1'b0;
assign w_ex1_rs2_mispred = r_ex1_issue.rd_regs[1].valid & r_ex1_issue.rd_regs[1].predict_ready ? w_ex1_rs2_lsu_mispred : 1'b0;

assign o_ex1_early_wr.valid = r_ex1_issue.valid & r_ex1_issue.wr_reg.valid &
                              ~w_ex1_rs1_mispred & ~w_ex1_rs2_mispred;
assign o_ex1_early_wr.rd_rnid = r_ex1_issue.wr_reg.rnid;
assign o_ex1_early_wr.rd_type = r_ex1_issue.wr_reg.typ;
assign o_ex1_early_wr.may_mispred = 1'b0;

generate
  for (genvar tgt_idx = 0; tgt_idx < msrh_pkg::REL_BUS_SIZE; tgt_idx++) begin : rs_tgt_loop
    assign w_ex2_rs1_fwd_valid[tgt_idx] = r_ex2_issue.rd_regs[0].valid & ex1_i_phy_wr[tgt_idx].valid &
                                          (r_ex2_issue.rd_regs[0].typ  == ex1_i_phy_wr[tgt_idx].rd_type) &
                                          (r_ex2_issue.rd_regs[0].rnid == ex1_i_phy_wr[tgt_idx].rd_rnid) &
                                          (r_ex2_issue.rd_regs[0].rnid != 'h0);   // GPR[x0] always zero

    assign w_ex2_rs2_fwd_valid[tgt_idx] = r_ex2_issue.rd_regs[1].valid & ex1_i_phy_wr[tgt_idx].valid &
                                          (r_ex2_issue.rd_regs[1].typ  == ex1_i_phy_wr[tgt_idx].rd_type) &
                                          (r_ex2_issue.rd_regs[1].rnid == ex1_i_phy_wr[tgt_idx].rd_rnid) &
                                          (r_ex2_issue.rd_regs[1].rnid != 'h0);   // GPR[x0] always zero
    assign w_ex2_tgt_data[tgt_idx] = ex1_i_phy_wr[tgt_idx].rd_data;
  end
endgenerate

bit_oh_or #(
    .T(riscv_pkg::xlen_t),
    .WORDS(msrh_pkg::TGT_BUS_SIZE)
) u_rs1_data_select (
    .i_oh(w_ex2_rs1_fwd_valid),
    .i_data(w_ex2_tgt_data),
    .o_selected(w_ex2_rs1_fwd_data)
);

bit_oh_or #(
    .T(riscv_pkg::xlen_t),
    .WORDS(msrh_pkg::TGT_BUS_SIZE)
) u_rs2_data_select (
    .i_oh(w_ex2_rs2_fwd_valid),
    .i_data(w_ex2_tgt_data),
    .o_selected(w_ex2_rs2_fwd_data)
);

// EX1 brtag flush check
assign w_ex1_br_flush  = msrh_pkg::is_br_flush_target(r_ex1_issue.br_mask, ex3_br_upd_if.brtag,
                                                      ex3_br_upd_if.dead, ex3_br_upd_if.mispredict) & ex3_br_upd_if.update & r_ex1_issue.valid;

always_comb begin
  w_ex2_issue_next = r_ex1_issue;
end

always_ff @(posedge i_clk, negedge i_reset_n) begin
  if (!i_reset_n) begin
    r_ex2_rs1_data <= 'h0;
    r_ex2_rs2_data <= 'h0;

    r_ex2_issue <= 'h0;
    r_ex2_index <= 'h0;
    r_ex2_pipe_ctrl <= 'h0;
    r_ex2_dead <= 1'b0;

    r_ex2_wr_valid <= 1'b0;
  end else begin
    r_ex2_rs1_data <= ex1_regread_rs1.data;
    r_ex2_rs2_data <= ex1_regread_rs2.data;

    r_ex2_issue <= w_ex2_issue_next;
    r_ex2_index <= r_ex1_index;
    r_ex2_pipe_ctrl <= r_ex1_pipe_ctrl;
    r_ex2_dead <= r_ex1_dead | r_ex1_issue.valid & (w_ex1_br_flush | w_commit_flushed);

    r_ex2_wr_valid <= o_ex1_early_wr.valid;
  end
end

assign w_ex2_rs1_selected_data = |w_ex2_rs1_fwd_valid ? w_ex2_rs1_fwd_data : r_ex2_rs1_data;
assign w_ex2_rs2_selected_data = |w_ex2_rs2_fwd_valid ? w_ex2_rs2_fwd_data : r_ex2_rs2_data;

assign w_ex2_rs1_pred_hit = r_ex2_issue.rd_regs[0].valid & r_ex2_issue.rd_regs[0].predict_ready ? |w_ex2_rs1_fwd_valid : 1'b1;
assign w_ex2_rs2_pred_hit = r_ex2_issue.rd_regs[1].valid & r_ex2_issue.rd_regs[1].predict_ready ? |w_ex2_rs2_fwd_valid : 1'b1;

// EX2 brtag flush check
assign w_ex2_br_flush  = msrh_pkg::is_br_flush_target(r_ex2_issue.br_mask, ex3_br_upd_if.brtag,
                                                      ex3_br_upd_if.dead, ex3_br_upd_if.mispredict) & ex3_br_upd_if.update & r_ex3_issue.valid;

always_comb begin
  w_ex3_issue_next = r_ex2_issue;
end

always_ff @(posedge i_clk, negedge i_reset_n) begin
  if (!i_reset_n) begin
    r_ex3_result   <= 'h0;
    r_ex3_index    <= 'h0;
    r_ex3_issue    <= 'h0;
    r_ex3_br_vaddr <= 'h0;
    r_ex3_pipe_ctrl <= 'h0;
    r_ex3_dead <= 1'b0;

    r_ex3_rs1_pred_hit <= 1'b0;
    r_ex3_rs2_pred_hit <= 1'b0;
  end else begin
    r_ex3_issue    <= w_ex3_issue_next;
    r_ex3_index    <= r_ex2_index;
    r_ex3_br_vaddr <= w_ex2_br_vaddr;
    r_ex3_pipe_ctrl <= r_ex2_pipe_ctrl;
    r_ex3_dead <= r_ex2_dead | r_ex2_issue.valid & (w_ex2_br_flush | w_commit_flushed);

    r_ex3_rs1_pred_hit <= w_ex2_rs1_pred_hit;
    r_ex3_rs2_pred_hit <= w_ex2_rs2_pred_hit;

    case (r_ex2_pipe_ctrl.op)
      OP_EQ : r_ex3_result <= w_ex2_rs1_selected_data == w_ex2_rs2_selected_data;
      OP_NE : r_ex3_result <= w_ex2_rs1_selected_data != w_ex2_rs2_selected_data;
      OP_LT : r_ex3_result <= $signed(w_ex2_rs1_selected_data) <  $signed(w_ex2_rs2_selected_data);
      OP_GE : r_ex3_result <= $signed(w_ex2_rs1_selected_data) >= $signed(w_ex2_rs2_selected_data);
      OP_LTU: r_ex3_result <= w_ex2_rs1_selected_data <  w_ex2_rs2_selected_data;
      OP_GEU: r_ex3_result <= w_ex2_rs1_selected_data >= w_ex2_rs2_selected_data;
      OP__  : r_ex3_result <= 1'b1;   // Unconditional Jump
      default : r_ex3_result <= 1'bx;
    endcase
  end
end

assign o_ex3_phy_wr.valid   = r_ex3_issue.valid &
                              r_ex3_pipe_ctrl.wr_rd & (r_ex3_issue.wr_reg.regidx != 'h0) &
                              r_ex3_rs1_pred_hit & r_ex3_rs2_pred_hit;
assign o_ex3_phy_wr.rd_rnid = r_ex3_issue.wr_reg.rnid;
assign o_ex3_phy_wr.rd_type = r_ex3_issue.wr_reg.typ;
assign o_ex3_phy_wr.rd_data = {{(riscv_pkg::XLEN_W-riscv_pkg::VADDR_W){r_ex3_issue.pc_addr[riscv_pkg::VADDR_W-1]}},
                               r_ex3_issue.pc_addr} + (r_ex3_issue.is_rvc ? 'h2 : 'h4);

assign ex3_done_if.done     = r_ex3_issue.valid & r_ex3_rs1_pred_hit & r_ex3_rs2_pred_hit;
assign ex3_done_if.index_oh = r_ex3_index;
assign ex3_done_if.except_valid  = 1'b0;
assign ex3_done_if.except_type = msrh_pkg::except_t'('h0);

logic [riscv_pkg::VADDR_W-1: 0] w_ex2_offset_uj;
logic [riscv_pkg::VADDR_W-1: 0] w_ex2_offset_sb;

assign w_ex2_offset_uj = {{(riscv_pkg::VADDR_W-21){r_ex2_issue.inst[31]}},
                          r_ex2_issue.inst[31],
                          r_ex2_issue.inst[19:12],
                          r_ex2_issue.inst[20],
                          r_ex2_issue.inst[30:21],
                          1'b0};
assign w_ex2_offset_sb = {{(riscv_pkg::VADDR_W-13){r_ex2_issue.inst[31]}},
                          r_ex2_issue.inst[31],
                          r_ex2_issue.inst[ 7],
                          r_ex2_issue.inst[30:25],
                          r_ex2_issue.inst[11: 8],
                          1'b0};

always_comb begin
  case (r_ex2_pipe_ctrl.imm)
    IMM_SB : w_ex2_br_vaddr = r_ex2_issue.pc_addr + w_ex2_offset_sb;
    IMM_UJ : w_ex2_br_vaddr = r_ex2_issue.pc_addr + w_ex2_offset_uj;
    IMM_I  : begin
      logic [riscv_pkg::VADDR_W-1: 0]          w_ex2_br_vaddr_tmp;
      w_ex2_br_vaddr_tmp = w_ex2_rs1_selected_data[riscv_pkg::VADDR_W-1: 0] +
                           {{(riscv_pkg::VADDR_W-12){r_ex2_issue.inst[31]}},
                            r_ex2_issue.inst[31:20]};
      // When JALR, clearing lowest bit
      w_ex2_br_vaddr = {w_ex2_br_vaddr_tmp[riscv_pkg::VADDR_W-1: 1], 1'b0};
    end
    default : w_ex2_br_vaddr = {riscv_pkg::VADDR_W{1'bx}};
  endcase // case (w_ex2_pipe_ctrl.imm)
end // always_comb

// logic w_ex3_not_predict_taken;
logic w_ex3_ras_hit;
logic w_ex3_bim_hit;

assign w_ex3_ras_hit = r_ex3_issue.is_ret & r_ex3_issue.pred_taken & (r_ex3_br_vaddr == r_ex3_issue.pred_target_vaddr);
assign w_ex3_bim_hit = r_ex3_issue.btb_valid &
                       ((~r_ex3_result & ~r_ex3_issue.pred_taken) |
                        (r_ex3_result & r_ex3_issue.pred_taken &
                         (r_ex3_br_vaddr == r_ex3_issue.pred_target_vaddr)));

assign ex3_br_upd_if.update        = r_ex3_issue.valid & r_ex3_rs1_pred_hit & r_ex3_rs2_pred_hit;
assign ex3_br_upd_if.is_call       = r_ex3_issue.is_call;
assign ex3_br_upd_if.is_ret        = r_ex3_issue.is_ret;
assign ex3_br_upd_if.is_rvc        = r_ex3_issue.is_rvc;
assign ex3_br_upd_if.ras_index     = r_ex3_issue.ras_index;
assign ex3_br_upd_if.taken         = r_ex3_result;
assign ex3_br_upd_if.dead          = r_ex3_dead;
assign ex3_br_upd_if.mispredict    = ~w_ex3_ras_hit & ~w_ex3_bim_hit;

assign ex3_br_upd_if.bim_value     = r_ex3_issue.bim_value;
assign ex3_br_upd_if.pc_vaddr      = /* r_ex3_issue.is_rvc ? */ r_ex3_issue.pc_addr /* : r_ex3_issue.pc_addr + 'h2 */;
assign ex3_br_upd_if.target_vaddr  = r_ex3_result ? r_ex3_br_vaddr :
                                     r_ex3_issue.is_rvc ? r_ex3_issue.pc_addr + 'h2 : r_ex3_issue.pc_addr + 'h4;
`ifdef SIMULATION
assign ex3_br_upd_if.pred_vaddr    = r_ex3_issue.pred_target_vaddr;
`endif // SIMULATION

assign ex3_br_upd_if.cmt_id        = r_ex3_issue.cmt_id;
assign ex3_br_upd_if.grp_id        = r_ex3_issue.grp_id;
assign ex3_br_upd_if.brtag         = r_ex3_issue.brtag;
assign ex3_br_upd_if.br_mask       = r_ex3_issue.br_mask;

`ifdef SIMULATION
`ifdef MONITOR

integer bim_fp;
initial begin
  bim_fp = $fopen("bru_detail.log", "w");
end

always_ff @ (negedge i_clk, negedge i_reset_n) begin
  if (i_reset_n) begin
    if (ex3_br_upd_if.update & ~ex3_br_upd_if.dead) begin
      if (r_ex3_pipe_ctrl.op != OP__) begin
        $fwrite(bim_fp, "%t : (%02d,%d) pc_vaddr = %08x, target_addr = %08x, %s, bim=%1d, %s, DASM(0x%08x)\n",
                $time,
                r_ex3_issue.cmt_id, r_ex3_issue.grp_id,
                r_ex3_issue.pc_addr,
                ex3_br_upd_if.target_vaddr,
                r_ex3_result ? "Taken   " : "NotTaken",
                ex3_br_upd_if.bim_value,
                ex3_br_upd_if.mispredict ? "Miss" : "Succ",
                r_ex3_issue.inst);
      end else if (r_ex3_issue.is_ret | r_ex3_issue.is_call) begin
        $fwrite(bim_fp, "%t : (%02d,%d) pc_vaddr = %08x, target_addr = %08x, pred_target_addr = %08x, ras_index = %d, %s, DASM(0x%08x)\n",
                $time,
                r_ex3_issue.cmt_id, r_ex3_issue.grp_id,
                r_ex3_issue.pc_addr,
                ex3_br_upd_if.target_vaddr,
                r_ex3_issue.pred_target_vaddr,
                r_ex3_issue.ras_index,
                ex3_br_upd_if.mispredict ? "Miss" : "Succ",
                r_ex3_issue.inst);
      end
    end
  end
  // if (msrh_tb.u_msrh_tile_wrapper.u_msrh_tile.u_frontend.u_predictor.u_ras.i_wr_valid) begin
  //   $fwrite(bim_fp, "%t : pc_vaddr = %08x, target_addr = %08x, pred_target_addr = %08x, ras_idx=%1d, %s, DASM(0x%08x)\n",
  //           $time,
  //           r_ex3_issue.pc_addr,
  //           ex3_br_upd_if.target_vaddr,
  //           r_ex3_issue.pred_target_vaddr,
  //           r_ex3_issue.ras_index,
  //           r_ex3_issue.inst);
  // end
end // always_ff @ (negedge i_clk, negedge i_reset_n)

final begin
  $fclose(bim_fp);
end

`endif // MONITOR
`endif // SIMULATION

endmodule // msrh_bru_pipe
