package riscv_common_pkg;

  // Privilege Mode
  localparam PRIV_U = 2'h0;
  localparam PRIV_S = 2'h1;
  localparam PRIV_H = 2'h2;
  localparam PRIV_M = 2'h3;

endpackage
