package riscv_fpu_pkg;

  localparam FLEN_W = 64;

endpackage // riscv_fpu_pkg
