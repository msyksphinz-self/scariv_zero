package msrh_fpu_pkg;

import decoder_fpu_ctrl_pkg::*;

endpackage // msrh_fpu_pkg
