riscv_fpu_imac_pkg.sv