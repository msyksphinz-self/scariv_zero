riscv_fpu_imfdc_pkg.sv