// ------------------------------------------------------------------------
// NAME : scariv_lsu_replay_queue
// TYPE : module
// ------------------------------------------------------------------------
// LSU Replay Queue
// ------------------------------------------------------------------------
//
// ------------------------------------------------------------------------

module scariv_lsu_replay_queue
  import scariv_lsu_pkg::*;
(
    input logic i_clk,
    input logic i_reset_n,

    input scariv_pkg::commit_blk_t i_commit,
    br_upd_if.slave                br_upd_if,

    lsu_pipe_haz_if.slave  lsu_pipe_haz_if,

    input missu_resolve_t  i_missu_resolve,
    input logic            i_missu_is_full,   

    // Request from Replay Queue
    lsu_pipe_req_if.master lsu_pipe_req_if
);

localparam REPLAY_QUEUE_SIZE = (scariv_conf_pkg::LDQ_SIZE + scariv_conf_pkg::STQ_SIZE) / 2;
localparam REPLAY_QUEUE_W = $clog2(REPLAY_QUEUE_SIZE);

logic [REPLAY_QUEUE_W-1: 0] r_diff_counter;

typedef struct packed {
    logic [31: 0]                                  inst;
    decoder_inst_cat_pkg::inst_cat_t               cat;
    logic                                          oldest_valid;
    scariv_pkg::reg_rd_issue_t                     rd_reg;
    scariv_pkg::reg_wr_issue_t                     wr_reg;
    scariv_pkg::paddr_t                            paddr;
    scariv_lsu_pkg::ex2_haz_t                      hazard_typ;
    logic [scariv_conf_pkg::MISSU_ENTRY_SIZE-1: 0] missu_index_oh;
    logic [REPLAY_QUEUE_W-1: 0]                    diff_counter;
} replay_queue_t;
typedef struct packed {
    logic                valid;
    logic                dead;
    scariv_pkg::cmt_id_t cmt_id;
    scariv_pkg::grp_id_t grp_id;
    scariv_pkg::brmask_t br_mask;
} replay_additional_queue_t;

replay_queue_t w_new_replay_queue_info;
replay_queue_t w_rd_replay_queue_info;
replay_additional_queue_t r_replay_additional_queue[REPLAY_QUEUE_SIZE];
logic w_lsu_replay_valid;

logic w_empty;
logic w_full;
logic w_queue_push;
logic w_queue_pop;

assign lsu_pipe_haz_if.full = w_full;
assign w_queue_push = lsu_pipe_haz_if.valid & !lsu_pipe_haz_if.full;
assign w_queue_pop  = w_lsu_replay_valid & lsu_pipe_req_if.ready;

assign w_new_replay_queue_info.inst           = lsu_pipe_haz_if.payload.inst          ;
assign w_new_replay_queue_info.cat            = lsu_pipe_haz_if.payload.cat           ;
assign w_new_replay_queue_info.oldest_valid   = lsu_pipe_haz_if.payload.oldest_valid  ;
assign w_new_replay_queue_info.rd_reg         = lsu_pipe_haz_if.payload.rd_reg        ;
assign w_new_replay_queue_info.wr_reg         = lsu_pipe_haz_if.payload.wr_reg        ;
assign w_new_replay_queue_info.paddr          = lsu_pipe_haz_if.payload.paddr         ;
assign w_new_replay_queue_info.hazard_typ     = lsu_pipe_haz_if.payload.hazard_typ    ;
assign w_new_replay_queue_info.missu_index_oh = lsu_pipe_haz_if.payload.missu_index_oh;
assign w_new_replay_queue_info.diff_counter   = r_diff_counter;

// Diff counter from previous Queue inesrtion
always_ff @ (posedge i_clk, negedge i_reset_n) begin
    if (!i_reset_n) begin
        r_diff_counter <= 'h0;
    end else begin
        if (w_empty) begin
            r_diff_counter <= 'h0;
        end else begin
            r_diff_counter <= r_diff_counter + 'h1;
        end
    end
end
logic [REPLAY_QUEUE_W-1: 0] r_replay_queue_head_ptr;
logic [REPLAY_QUEUE_W-1: 0] r_replay_queue_tail_ptr;
generate for (genvar idx = 0; idx < REPLAY_QUEUE_SIZE; idx++) begin : replay_additional_loop
    logic w_commit_flush;
    logic w_br_flush;
    logic w_entry_flush;
    assign w_commit_flush = scariv_pkg::is_commit_flush_target(r_replay_additional_queue[idx].cmt_id, 
                                                               r_replay_additional_queue[idx].grp_id, 
                                                               i_commit) & r_replay_additional_queue[idx].valid;
    assign w_br_flush     = scariv_pkg::is_br_flush_target(r_replay_additional_queue[idx].br_mask, br_upd_if.brtag,
                                                           br_upd_if.dead, br_upd_if.mispredict) & br_upd_if.update & r_replay_additional_queue[idx].valid;
    assign w_entry_flush  = w_commit_flush | w_br_flush;

    always_ff @ (posedge i_clk, negedge i_reset_n) begin
        if (w_queue_push & 
            (idx == r_replay_queue_head_ptr)) begin
            r_replay_additional_queue[idx].valid   <= 1'b1;
            r_replay_additional_queue[idx].dead    <= 1'b0;
            r_replay_additional_queue[idx].cmt_id  <= lsu_pipe_haz_if.payload.cmt_id;
            r_replay_additional_queue[idx].grp_id  <= lsu_pipe_haz_if.payload.grp_id;
            r_replay_additional_queue[idx].br_mask <= lsu_pipe_haz_if.payload.br_mask;
        end else if (w_queue_pop &
                (idx == r_replay_queue_tail_ptr)) begin
            r_replay_additional_queue[idx].valid  <= 1'b0;
        end else if (r_replay_additional_queue[idx].valid &
                     w_entry_flush) begin
            r_replay_additional_queue[idx].dead <= 1'b1;
        end
    end
end endgenerate

always_ff @ (posedge i_clk, negedge i_reset_n) begin
    if (!i_reset_n) begin
        r_replay_queue_head_ptr <= 'h0;
        r_replay_queue_tail_ptr <= 'h0;        
    end else begin
        if (w_queue_push) begin
            r_replay_queue_head_ptr <= r_replay_queue_head_ptr + 'h1;
        end
        if (w_queue_pop) begin
            r_replay_queue_tail_ptr <= r_replay_queue_tail_ptr + 'h1;
        end
    end
end

ring_fifo
#(
    .T     (replay_queue_t),
    .DEPTH (REPLAY_QUEUE_SIZE)
)
u_replay_queue
(
    .i_clk     (i_clk    ),
    .i_reset_n (i_reset_n),

    .i_push (w_queue_push  ),
    .i_data (w_new_replay_queue_info),

    .o_empty(w_empty),
    .o_full (w_full ),

    .i_pop  (w_queue_pop),
    .o_data (w_rd_replay_queue_info)
);

logic [REPLAY_QUEUE_W-1: 0] r_prev_diff_counter;

always_ff @ (posedge i_clk, negedge i_reset_n) begin
    if (!i_reset_n) begin
        r_prev_diff_counter <= 'h0;
    end else begin
        if (w_queue_pop) begin
            r_prev_diff_counter <= 'h0;
        end else begin
            r_prev_diff_counter <= r_prev_diff_counter + 'h1;
        end
    end
end

always_comb begin
    if (!w_empty) begin
        if (w_rd_replay_queue_info.diff_counter != 'h0 && 
            r_prev_diff_counter == w_rd_replay_queue_info.diff_counter) begin
            w_lsu_replay_valid = !r_replay_additional_queue[r_replay_queue_tail_ptr].dead;
        end else begin
            case (w_rd_replay_queue_info.hazard_typ)
                EX2_HAZ_STQ_NONFWD_HAZ : w_lsu_replay_valid = 1'b0; 
                EX2_HAZ_RMW_ORDER_HAZ :  w_lsu_replay_valid = 1'b0;
                EX2_HAZ_L1D_CONFLICT :   w_lsu_replay_valid = 1'b1; // Replay immediately
                EX2_HAZ_MISSU_FULL :     w_lsu_replay_valid = i_missu_is_full;
                EX2_HAZ_MISSU_ASSIGNED : w_lsu_replay_valid = i_missu_resolve.valid & (i_missu_resolve.resolve_index_oh == w_rd_replay_queue_info.missu_index_oh);
                default : begin
                    w_lsu_replay_valid = 1'b0;
                    // $fatal(0, "Must not come here. hazard_typ = %d", w_rd_replay_queue_info.hazard_typ);
                end
            endcase
        end
    end else begin
        w_lsu_replay_valid = 1'b0;
    end

    lsu_pipe_req_if.payload.cmt_id         = r_replay_additional_queue[r_replay_queue_tail_ptr].cmt_id;
    lsu_pipe_req_if.payload.grp_id         = r_replay_additional_queue[r_replay_queue_tail_ptr].grp_id;
    lsu_pipe_req_if.payload.br_mask        = r_replay_additional_queue[r_replay_queue_tail_ptr].br_mask;
    lsu_pipe_req_if.payload.inst           = w_rd_replay_queue_info.inst          ;
    lsu_pipe_req_if.payload.cat            = w_rd_replay_queue_info.cat           ;
    lsu_pipe_req_if.payload.oldest_valid   = w_rd_replay_queue_info.oldest_valid  ;
    lsu_pipe_req_if.payload.rd_reg         = w_rd_replay_queue_info.rd_reg        ;
    lsu_pipe_req_if.payload.wr_reg         = w_rd_replay_queue_info.wr_reg        ;
    lsu_pipe_req_if.payload.paddr          = w_rd_replay_queue_info.paddr         ;
    lsu_pipe_req_if.payload.hazard_typ     = w_rd_replay_queue_info.hazard_typ    ;
    lsu_pipe_req_if.payload.missu_index_oh = w_rd_replay_queue_info.missu_index_oh;
    
end
assign lsu_pipe_req_if.valid = w_lsu_replay_valid & ~r_replay_additional_queue[r_replay_queue_tail_ptr].dead;

`ifdef SIMULATION
always_ff @ (negedge i_clk, negedge i_reset_n) begin
    if (i_reset_n) begin
        if (!w_empty) begin
            case (w_rd_replay_queue_info.hazard_typ)
                EX2_HAZ_STQ_NONFWD_HAZ : begin end  
                EX2_HAZ_RMW_ORDER_HAZ :  begin end 
                EX2_HAZ_L1D_CONFLICT :   begin end
                EX2_HAZ_MISSU_FULL :     begin end
                EX2_HAZ_MISSU_ASSIGNED : begin end
                default : begin
                    $fatal(0, "Must not come here. hazard_typ = %d", w_rd_replay_queue_info.hazard_typ);
                end
            endcase
        end
    end
end
`endif // SIMULATION


endmodule
