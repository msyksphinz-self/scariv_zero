`define RV64
