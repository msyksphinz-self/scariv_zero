module msrh_bru_rn_snapshots    //
  import msrh_pkg::*;
  (
   input logic         i_clk,
   input logic         i_reset_n,

   input rnid_t i_rn_list[32],

   input grp_id_t      i_load,
   input grp_id_t      i_rd_valid,
   input logic [ 4: 0] i_rd_archreg[msrh_conf_pkg::DISP_SIZE],
   input rnid_t        i_rd_rnid   [msrh_conf_pkg::DISP_SIZE],
   input brtag_t       i_brtag     [msrh_conf_pkg::DISP_SIZE],

   // Branch Tag Update Signal
   br_upd_if.slave br_upd_if,

   output              rnid_t o_rn_list[32]
   );

logic [31: 0][RNID_W-1: 0] r_snapshots[msrh_conf_pkg::RV_BRU_ENTRY_SIZE];
/* verilator lint_off UNOPTFLAT */
logic [31: 0][RNID_W-1: 0] w_tmp_snapshots[msrh_conf_pkg::DISP_SIZE+1];

generate for(genvar i =  0; i < 32; i++) begin
  assign w_tmp_snapshots[0][i] = i_rn_list[i];
end
endgenerate

brtag_t w_brtag_sel;
bit_oh_or #(.T(brtag_t), .WORDS(msrh_conf_pkg::DISP_SIZE))
u_brtag_sel (.i_oh(i_load), .i_data(i_brtag), .o_selected(w_brtag_sel));


generate for(genvar r_idx =  0; r_idx < 32; r_idx++) begin : register_loop
  for (genvar d_idx = 0; d_idx < msrh_conf_pkg::DISP_SIZE; d_idx++) begin : disp_loop
    /* verilator lint_off ALWCOMBORDER */
    assign w_tmp_snapshots[d_idx+1][r_idx] = i_rd_valid[d_idx] & (i_rd_archreg[d_idx] == r_idx[ 4: 0]) ? i_rd_rnid[d_idx] : w_tmp_snapshots[d_idx][r_idx[ 4: 0]];
  end

end
endgenerate

generate for (genvar i_idx = 0; i_idx < 32; i_idx++) begin : reg_loop
  always_ff @ (posedge i_clk) begin
    if (|i_load) begin
      r_snapshots[i_brtag[0]][i_idx] <= w_tmp_snapshots[msrh_conf_pkg::DISP_SIZE][i_idx];
    end
  end
end
endgenerate

generate for(genvar i =  0; i < 32; i++) begin : o_loop
  assign o_rn_list[i] = r_snapshots[br_upd_if.brtag][i];
end
endgenerate

endmodule // msrh_bru_rn_snapshots
