riscv_fpu_imc_pkg.sv