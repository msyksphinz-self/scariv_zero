kimura@kimura-tower.3065934:1708515676