module msrh_ras
  (
   input logic                                              i_clk,
   input logic                                              i_reset,

   input logic                                              i_wr_valid,
   input logic [$clog2(msrh_conf_pkg::RAS_ENTRY_SIZE)-1:0]  i_wr_index,
   input logic [riscv_pkg::PADDR_W-1: 0]                    i_wr_pa,

   output logic                                             i_rd_valid,
   output logic [$clog2(msrh_conf_pkg::RAS_ENTRY_SIZE)-1:0] i_rd_index,
   output logic [riscv_pkg::PADDR_W-1: 0]                   o_rd_pa
   );

logic [PADDR_W-1: 0] r_ras_array[msrh_conf_pkg::RAS_ENTRY_SIZE];

always_ff @ (posedge i_clk, negedge i_reset_n) begin
  if (!i_reset_n) begin
    for (int i = 0; i < msrh_conf_pkg::RAS_ENTRY_SIZE; i++) begin
      r_ras_array[i] <= 'h0;
    end
  end else begin
    if (i_wr_valid) begin
      r_ras_array[i_wr_index] <= i_wr_pa;
    end
  end
end

assign o_rd_pa = i_rd_valid ? r_ras_array[i_rd_index] : 'h0;

endmodule // msrh_ras
