package riscv_common_pkg;

  // Privilege Mode
  localparam RRIV_U = 2'h0;
  localparam RRIV_S = 2'h1;
  localparam RRIV_H = 2'h2;
  localparam RRIV_M = 2'h3;

endpackage
