package msrh_conf_pkg;

  localparam DISP_SIZE = 3;

  localparam ALU_INST_NUM = 1;
  localparam LSU_INST_NUM = 1;

  localparam ARITH_DISP_SIZE = 2;
  localparam MEM_DISP_SIZE = 2;

endpackage // msrh_conf_pkg
