package riscv_fpu_pkg;

  localparam FLEN_W = 32;

endpackage // riscv_fpu_pkg
