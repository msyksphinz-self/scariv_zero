`define RV64
`define LITEX_SIMULATION
`define RV_AMO 1
