`define SYSREG_ADDR_USTATUS 12'h000
`define SYSREG_ADDR_UIE 12'h004
`define SYSREG_ADDR_UTVEC 12'h005
`define SYSREG_ADDR_VSTART 12'h008
`define SYSREG_ADDR_VXSAT 12'h009
`define SYSREG_ADDR_VXRM 12'h00a
`define SYSREG_ADDR_USCRATCH 12'h040
`define SYSREG_ADDR_UEPC 12'h041
`define SYSREG_ADDR_UCAUSE 12'h042
`define SYSREG_ADDR_UBADADDR 12'h043
`define SYSREG_ADDR_UIP 12'h044
`define SYSREG_ADDR_FFLAGS 12'h001
`define SYSREG_ADDR_FRM 12'h002
`define SYSREG_ADDR_FCSR 12'h003
`define SYSREG_ADDR_CYCLE 12'hc00
`define SYSREG_ADDR_TIME  12'hc01
`define SYSREG_ADDR_INSTRET 12'hc02
`define SYSREG_ADDR_HPMCOUNTER3 12'hc03
`define SYSREG_ADDR_HPMCOUNTER4 12'hc04
`define SYSREG_ADDR_HPMCOUNTER5 12'hc05
`define SYSREG_ADDR_HPMCOUNTER6 12'hc06
`define SYSREG_ADDR_HPMCOUNTER7 12'hc07
`define SYSREG_ADDR_HPMCOUNTER8 12'hc08
`define SYSREG_ADDR_HPMCOUNTER9 12'hc09
`define SYSREG_ADDR_HPMCOUNTER10 12'hc0a
`define SYSREG_ADDR_HPMCOUNTER11 12'hc0b
`define SYSREG_ADDR_HPMCOUNTER12 12'hc0c
`define SYSREG_ADDR_HPMCOUNTER13 12'hc0d
`define SYSREG_ADDR_HPMCOUNTER14 12'hc0e
`define SYSREG_ADDR_HPMCOUNTER15 12'hc0f
`define SYSREG_ADDR_HPMCOUNTER16 12'hc10
`define SYSREG_ADDR_HPMCOUNTER17 12'hc11
`define SYSREG_ADDR_HPMCOUNTER18 12'hc12
`define SYSREG_ADDR_HPMCOUNTER19 12'hc13
`define SYSREG_ADDR_HPMCOUNTER20 12'hc14
`define SYSREG_ADDR_HPMCOUNTER21 12'hc15
`define SYSREG_ADDR_HPMCOUNTER22 12'hc16
`define SYSREG_ADDR_HPMCOUNTER23 12'hc17
`define SYSREG_ADDR_HPMCOUNTER24 12'hc18
`define SYSREG_ADDR_HPMCOUNTER25 12'hc19
`define SYSREG_ADDR_HPMCOUNTER26 12'hc1a
`define SYSREG_ADDR_HPMCOUNTER27 12'hc1b
`define SYSREG_ADDR_HPMCOUNTER28 12'hc1c
`define SYSREG_ADDR_HPMCOUNTER29 12'hc1d
`define SYSREG_ADDR_HPMCOUNTER30 12'hc1e
`define SYSREG_ADDR_HPMCOUNTER31 12'hc1f
`define SYSREG_ADDR_CYCLEH 12'hc80
`define SYSREG_ADDR_TIMEH 12'hc81
`define SYSREG_ADDR_INSTRETH 12'hc82
`define SYSREG_ADDR_HPMCOUNTERH3 12'hc83
`define SYSREG_ADDR_HPMCOUNTERH4 12'hc84
`define SYSREG_ADDR_HPMCOUNTERH5 12'hc85
`define SYSREG_ADDR_HPMCOUNTERH6 12'hc86
`define SYSREG_ADDR_HPMCOUNTERH7 12'hc87
`define SYSREG_ADDR_HPMCOUNTERH8 12'hc88
`define SYSREG_ADDR_HPMCOUNTERH9 12'hc89
`define SYSREG_ADDR_HPMCOUNTERH10 12'hc8a
`define SYSREG_ADDR_HPMCOUNTERH11 12'hc8b
`define SYSREG_ADDR_HPMCOUNTERH12 12'hc8c
`define SYSREG_ADDR_HPMCOUNTERH13 12'hc8d
`define SYSREG_ADDR_HPMCOUNTERH14 12'hc8e
`define SYSREG_ADDR_HPMCOUNTERH15 12'hc8f
`define SYSREG_ADDR_HPMCOUNTERH16 12'hc90
`define SYSREG_ADDR_HPMCOUNTERH17 12'hc91
`define SYSREG_ADDR_HPMCOUNTERH18 12'hc92
`define SYSREG_ADDR_HPMCOUNTERH19 12'hc93
`define SYSREG_ADDR_HPMCOUNTERH20 12'hc94
`define SYSREG_ADDR_HPMCOUNTERH21 12'hc95
`define SYSREG_ADDR_HPMCOUNTERH22 12'hc96
`define SYSREG_ADDR_HPMCOUNTERH23 12'hc97
`define SYSREG_ADDR_HPMCOUNTERH24 12'hc98
`define SYSREG_ADDR_HPMCOUNTERH25 12'hc99
`define SYSREG_ADDR_HPMCOUNTERH26 12'hc9a
`define SYSREG_ADDR_HPMCOUNTERH27 12'hc9b
`define SYSREG_ADDR_HPMCOUNTERH28 12'hc9c
`define SYSREG_ADDR_HPMCOUNTERH29 12'hc9d
`define SYSREG_ADDR_HPMCOUNTERH30 12'hc9e
`define SYSREG_ADDR_HPMCOUNTERH31 12'hc9f
`define SYSREG_ADDR_SSTATUS 12'h100
`define SYSREG_ADDR_SEDELEG 12'h102
`define SYSREG_ADDR_SIDELEG 12'h103
`define SYSREG_ADDR_SIE 12'h104
`define SYSREG_ADDR_STVEC 12'h105
`define SYSREG_ADDR_SCOUNTEREN 12'h106
`define SYSREG_ADDR_SSCRATCH 12'h140
`define SYSREG_ADDR_SEPC 12'h141
`define SYSREG_ADDR_SCAUSE 12'h142
`define SYSREG_ADDR_STVAL 12'h143
`define SYSREG_ADDR_SIP 12'h144
`define SYSREG_ADDR_SATP 12'h180
`define SYSREG_ADDR_HSTATUS 12'h200
`define SYSREG_ADDR_HEDELEG 12'h202
`define SYSREG_ADDR_HIDELEG 12'h203
`define SYSREG_ADDR_HIE 12'h204
`define SYSREG_ADDR_HTVEC 12'h205
`define SYSREG_ADDR_HSCRATCH 12'h240
`define SYSREG_ADDR_HEPC 12'h241
`define SYSREG_ADDR_HCAUSE 12'h242
`define SYSREG_ADDR_HBADADDR 12'h243
`define SYSREG_ADDR_HIP 12'h244
`define SYSREG_ADDR_HPTBR 12'h280
`define SYSREG_ADDR_MVENDORID 12'hf11
`define SYSREG_ADDR_MARCHID 12'hf12
`define SYSREG_ADDR_MIMPID 12'hf13
`define SYSREG_ADDR_MHARTID 12'hf14
`define SYSREG_ADDR_MSTATUS 12'h300
`define SYSREG_ADDR_MISA 12'h301
`define SYSREG_ADDR_MEDELEG 12'h302
`define SYSREG_ADDR_MIDELEG 12'h303
`define SYSREG_ADDR_MIE 12'h304
`define SYSREG_ADDR_MTVEC 12'h305
`define SYSREG_ADDR_MCOUNTEREN 12'h306
`define SYSREG_ADDR_MSCRATCH 12'h340
`define SYSREG_ADDR_MEPC 12'h341
`define SYSREG_ADDR_MCAUSE 12'h342
`define SYSREG_ADDR_MTVAL 12'h343
`define SYSREG_ADDR_MIP 12'h344
`define SYSREG_ADDR_MBASE 12'h380
`define SYSREG_ADDR_MBOUND 12'h381
`define SYSREG_ADDR_MIBASE 12'h382
`define SYSREG_ADDR_MIBOUND 12'h383
`define SYSREG_ADDR_MDBASE 12'h384
`define SYSREG_ADDR_MDBOUND 12'h385
`define SYSREG_ADDR_MCYCLE 12'hb00
`define SYSREG_ADDR_MINSTRET 12'hb02
`define SYSREG_ADDR_MHPMCOUNTER3 12'hb03
`define SYSREG_ADDR_MHPMCOUNTER4 12'hb04
`define SYSREG_ADDR_MHPMCOUNTER5 12'hb05
`define SYSREG_ADDR_MHPMCOUNTER6 12'hb06
`define SYSREG_ADDR_MHPMCOUNTER7 12'hb07
`define SYSREG_ADDR_MHPMCOUNTER8 12'hb08
`define SYSREG_ADDR_MHPMCOUNTER9 12'hb09
`define SYSREG_ADDR_MHPMCOUNTER10 12'hb0a
`define SYSREG_ADDR_MHPMCOUNTER11 12'hb0b
`define SYSREG_ADDR_MHPMCOUNTER12 12'hb0c
`define SYSREG_ADDR_MHPMCOUNTER13 12'hb0d
`define SYSREG_ADDR_MHPMCOUNTER14 12'hb0e
`define SYSREG_ADDR_MHPMCOUNTER15 12'hb0f
`define SYSREG_ADDR_MHPMCOUNTER16 12'hb10
`define SYSREG_ADDR_MHPMCOUNTER17 12'hb11
`define SYSREG_ADDR_MHPMCOUNTER18 12'hb12
`define SYSREG_ADDR_MHPMCOUNTER19 12'hb13
`define SYSREG_ADDR_MHPMCOUNTER20 12'hb14
`define SYSREG_ADDR_MHPMCOUNTER21 12'hb15
`define SYSREG_ADDR_MHPMCOUNTER22 12'hb16
`define SYSREG_ADDR_MHPMCOUNTER23 12'hb17
`define SYSREG_ADDR_MHPMCOUNTER24 12'hb18
`define SYSREG_ADDR_MHPMCOUNTER25 12'hb19
`define SYSREG_ADDR_MHPMCOUNTER26 12'hb1a
`define SYSREG_ADDR_MHPMCOUNTER27 12'hb1b
`define SYSREG_ADDR_MHPMCOUNTER28 12'hb1c
`define SYSREG_ADDR_MHPMCOUNTER29 12'hb1d
`define SYSREG_ADDR_MHPMCOUNTER30 12'hb1e
`define SYSREG_ADDR_MHPMCOUNTER31 12'hb1f
`define SYSREG_ADDR_MHPEVENT3 12'h323
`define SYSREG_ADDR_MHPEVENT4 12'h324
`define SYSREG_ADDR_MHPEVENT5 12'h325
`define SYSREG_ADDR_MHPEVENT6 12'h326
`define SYSREG_ADDR_MHPEVENT7 12'h327
`define SYSREG_ADDR_MHPEVENT8 12'h328
`define SYSREG_ADDR_MHPEVENT9 12'h329
`define SYSREG_ADDR_MHPEVENT10 12'h32a
`define SYSREG_ADDR_MHPEVENT11 12'h32b
`define SYSREG_ADDR_MHPEVENT12 12'h32c
`define SYSREG_ADDR_MHPEVENT13 12'h32d
`define SYSREG_ADDR_MHPEVENT14 12'h32e
`define SYSREG_ADDR_MHPEVENT15 12'h32f
`define SYSREG_ADDR_MHPEVENT16 12'h330
`define SYSREG_ADDR_MHPEVENT17 12'h331
`define SYSREG_ADDR_MHPEVENT18 12'h332
`define SYSREG_ADDR_MHPEVENT19 12'h333
`define SYSREG_ADDR_MHPEVENT20 12'h334
`define SYSREG_ADDR_MHPEVENT21 12'h335
`define SYSREG_ADDR_MHPEVENT22 12'h336
`define SYSREG_ADDR_MHPEVENT23 12'h337
`define SYSREG_ADDR_MHPEVENT24 12'h338
`define SYSREG_ADDR_MHPEVENT25 12'h339
`define SYSREG_ADDR_MHPEVENT26 12'h33a
`define SYSREG_ADDR_MHPEVENT27 12'h33b
`define SYSREG_ADDR_MHPEVENT28 12'h33c
`define SYSREG_ADDR_MHPEVENT29 12'h33d
`define SYSREG_ADDR_MHPEVENT30 12'h33e
`define SYSREG_ADDR_MHPEVENT31 12'h33f
`define SYSREG_ADDR_PMPCFG0 12'h3a0
`define SYSREG_ADDR_PMPCFG1 12'h3a1
`define SYSREG_ADDR_PMPCFG2 12'h3a2
`define SYSREG_ADDR_PMPCFG3 12'h3a3
`define SYSREG_ADDR_PMPADDR0 12'h3b0
`define SYSREG_ADDR_PMPADDR1 12'h3b1
`define SYSREG_ADDR_PMPADDR2 12'h3b2
`define SYSREG_ADDR_PMPADDR3 12'h3b3
`define SYSREG_ADDR_PMPADDR4 12'h3b4
`define SYSREG_ADDR_PMPADDR5 12'h3b5
`define SYSREG_ADDR_PMPADDR6 12'h3b6
`define SYSREG_ADDR_PMPADDR7 12'h3b7
`define SYSREG_ADDR_PMPADDR8 12'h3b8
`define SYSREG_ADDR_PMPADDR9 12'h3b9
`define SYSREG_ADDR_PMPADDR10 12'h3ba
`define SYSREG_ADDR_PMPADDR11 12'h3bb
`define SYSREG_ADDR_PMPADDR12 12'h3bc
`define SYSREG_ADDR_PMPADDR13 12'h3bd
`define SYSREG_ADDR_PMPADDR14 12'h3be
`define SYSREG_ADDR_PMPADDR15 12'h3bf
`define SYSREG_ADDR_STATS 12'h0c0

`define SYSREG_ADDR_SCONTEXT      12'h5a8
`define SYSREG_ADDR_TSELECT       12'h7a0
`define SYSREG_ADDR_TDATA1        12'h7a1
// `define SYSREG_ADDR_MCONTROL      12'h7a1
// `define SYSREG_ADDR_MCONTROL6     12'h7a1
// `define SYSREG_ADDR_ICOUNT        12'h7a1
// `define SYSREG_ADDR_ITRIGGER      12'h7a1
// `define SYSREG_ADDR_ETRIGGER      12'h7a1
// `define SYSREG_ADDR_TMEXTTRIGGER  12'h7a1
`define SYSREG_ADDR_TDATA2        12'h7a2
`define SYSREG_ADDR_TDATA3        12'h7a3
// `define SYSREG_ADDR_TEXT          12'h7a3
`define SYSREG_ADDR_TINFO         12'h7a4
`define SYSREG_ADDR_TCONTROL      12'h7a5
`define SYSREG_ADDR_MCONTEXT      12'h7a8
`define SYSREG_ADDR_MSCONTEXT     12'h7aa

`define MSTATUS_SIE  1
`define MSTATUS_SPIE 5
`define MSTATUS_SPP  8

`define MSTATUS_MIE  3
`define MSTATUS_MPIE 7
`define MSTATUS_MPP  12:11
`define MSTATUS_FS   14:13
`define MSTATUS_XS   16:15
`define MSTATUS_MPRV 17

`define MSTATUS_SUM 18
`define MSTATUS_MXR 19
`define MSTATUS_TVM 20
`define MSTATUS_TW  21
`define MSTATUS_TSR 22

`define SSTATUS_SIE  1
`define SSTATUS_SPIE 5
`define SSTATUS_SPP  8
