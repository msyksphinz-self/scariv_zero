`define RV64
`define RV_AMO (1)
// `define SIMULATION
// `define SUBSYSTEM_TOP sim.scariv_subsystem_axi_wrapper.u_scariv_subsystem
// `define NATIVE_DUMP
`define LITEX_FPGA
`define ILA_DEBUG
