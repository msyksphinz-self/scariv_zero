package msrh_conf_pkg;

  localparam DISP_SIZE = 8;

  localparam ALU_INST_NUM = 4;
  localparam LSU_INST_NUM = 3;

  localparam ARITH_DISP_SIZE = 8;
  localparam MEM_DISP_SIZE = 6;

endpackage // msrh_conf_pkg
