package sim_pkg;

localparam COUNT_UNIT = 1000;

endpackage // sim_pkg
