module select_early_wr_bus
  #(parameter REG_TYPE = scariv_pkg::GPR,
    localparam REN_UPD_NUM = REG_TYPE == scariv_pkg::GPR ? scariv_pkg::REL_XPR_BUS_SIZE : scariv_pkg::REL_FPR_BUS_SIZE
    )
(
   input scariv_pkg::rnid_t       i_entry_rnid,
   input scariv_pkg::reg_t        i_entry_type,
   input scariv_pkg::early_wr_t   i_early_wr[REN_UPD_NUM],

   output logic                 o_valid,
   output logic                 o_may_mispred
   );

logic [REN_UPD_NUM-1:0] w_rel_hit;
logic [REN_UPD_NUM-1:0] w_rel_hit_may_mispred;

scariv_pkg::early_wr_t alu_idx0, alu_idx1;
assign alu_idx0 = i_early_wr[0];
assign alu_idx1 = i_early_wr[1];


generate for (genvar r_idx = 0; r_idx < REN_UPD_NUM; r_idx++) begin : early_wr_loop
  assign w_rel_hit[r_idx] = i_early_wr[r_idx].valid &&
                            ((REG_TYPE == scariv_pkg::GPR) ? (i_early_wr[r_idx].rd_rnid != 'h0) : 1'b1) &
                            (i_entry_rnid == i_early_wr[r_idx].rd_rnid);
  assign w_rel_hit_may_mispred[r_idx] = w_rel_hit[r_idx] & i_early_wr[r_idx].may_mispred;
end endgenerate

assign o_valid = |w_rel_hit;
assign o_may_mispred = |w_rel_hit_may_mispred;

endmodule // select_early_wr_bus
