package riscv_vec_conf_pkg;

  parameter VLEN_W = 64;
  parameter DLEN_W = 64;

endpackage // riscv_vec_conf_pkg
