package riscv_vec_conf_pkg;

  parameter VLEN_W = 512;
  parameter DLEN_W = 128;

endpackage // riscv_vec_pkg
