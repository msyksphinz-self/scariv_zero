package riscv_vec_conf_pkg;

  parameter VLEN_W = 128;
  parameter DLEN_W = 128;

endpackage // riscv_vec_conf_pkg
