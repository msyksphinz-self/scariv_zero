package riscv_fpu_pkg;

  localparam FLEN_W = 0;

endpackage // riscv_fpu_pkg
