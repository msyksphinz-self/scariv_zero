module msrh_stq
  (
   );

endmodule // msrh_stq
