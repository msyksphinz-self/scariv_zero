package riscv_fpu_pkg;

parameter FLEN_W = 32;

endpackage // riscv_fpu_pkg
