module msrh_ldq
  import msrh_lsu_pkg::*;
(
   input logic                           i_clk,
   input logic                           i_reset_n,

   input logic [msrh_pkg::DISP_SIZE-1:0] i_disp_valid,
   disp_if.slave disp,

   // Updates from LSU Pipeline EX1 stage
   input ex1_q_update_t        i_ex1_q_updates[msrh_pkg::LSU_INST_NUM],
   // Updates from LSU Pipeline EX2 stage
   input logic [msrh_pkg::LSU_INST_NUM-1: 0] i_tlb_resolve,
   input ex2_q_update_t        i_ex2_q_updates[msrh_pkg::LSU_INST_NUM],

   lsu_replay_if.master ldq_replay_if[msrh_pkg::LSU_INST_NUM],

   input lrq_resolve_t     i_lrq_resolve,

   input logic [msrh_pkg::LSU_INST_NUM-1: 0] i_ex3_done,

   output                                msrh_pkg::done_rpt_t o_done_report
   );

ldq_entry_t w_ldq_entries[LDQ_SIZE];

msrh_pkg::disp_t disp_picked_inst[msrh_conf_pkg::MEM_DISP_SIZE];
logic [msrh_conf_pkg::MEM_DISP_SIZE-1:0] disp_picked_inst_valid;
logic [msrh_pkg::DISP_SIZE-1:0] disp_picked_grp_id[msrh_conf_pkg::MEM_DISP_SIZE];

logic [LDQ_SIZE-1: 0] w_rerun_request[msrh_pkg::LSU_INST_NUM];
logic [LDQ_SIZE-1: 0] w_rerun_request_oh[msrh_pkg::LSU_INST_NUM];
logic [msrh_pkg::LSU_INST_NUM-1: 0] w_rerun_request_rev_oh[LDQ_SIZE] ;
logic [msrh_pkg::LSU_INST_NUM-1: 0] w_ldq_replay_conflict[LDQ_SIZE] ;

//
// Done Selection
//
ldq_entry_t w_ldq_done_entry;
logic [LDQ_SIZE-1:0]  w_ldq_done_oh;

msrh_disp_pickup
  #(
    .PORT_BASE(0),
    .PORT_SIZE(msrh_conf_pkg::MEM_DISP_SIZE)
    )
u_msrh_disp_pickup
  (
   .i_disp_valid (i_disp_valid),
   .i_disp (disp),

   .o_disp_valid  (disp_picked_inst_valid),
   .o_disp        (disp_picked_inst),
   .o_disp_grp_id (disp_picked_grp_id)
   );

//
// LDQ Pointer
//
logic [$clog2(LDQ_SIZE)-1:0] w_in_ptr;
logic [$clog2(LDQ_SIZE)-1:0] w_out_ptr;
logic                                        w_in_vld;
logic                                        w_out_vld;
logic [LDQ_SIZE-1:0]         w_load_valid;
logic [$clog2(LDQ_SIZE):0]   w_disp_picked_num;

assign w_in_vld  = |disp_picked_inst_valid;
assign w_out_vld = o_done_report.valid;

/* verilator lint_off WIDTH */
bit_cnt #(.WIDTH(LDQ_SIZE)) cnt_disp_vld(.in({{(LDQ_SIZE-msrh_conf_pkg::MEM_DISP_SIZE){1'b0}}, disp_picked_inst_valid}), .out(w_disp_picked_num));
inoutptr_var #(.SIZE(LDQ_SIZE)) u_req_ptr(.i_clk (i_clk), .i_reset_n(i_reset_n),
                                                        .i_in_vld (w_in_vld ), .i_in_val (w_disp_picked_num[$clog2(LDQ_SIZE)-1: 0]), .o_in_ptr (w_in_ptr ),
                                                        .i_out_vld(w_out_vld), .i_out_val({{($clog2(LDQ_SIZE)-1){1'b0}}, 1'b1}), .o_out_ptr(w_out_ptr));

`ifdef SIMULATION
always_ff @ (negedge i_clk, negedge i_reset_n) begin
  if (!i_reset_n) begin
  end else begin
    if (w_disp_picked_num[$clog2(LDQ_SIZE)]) begin
      $fatal("w_disp_picked_num MSB == 1, too much requests inserted\n");
    end
  end
end
`endif // SIMULATION

generate for (genvar l_idx = 0; l_idx < LDQ_SIZE; l_idx++) begin : ldq_loop
  logic [msrh_conf_pkg::MEM_DISP_SIZE-1: 0]  w_input_valid;
  msrh_pkg::disp_t           w_disp_entry;
  logic [msrh_pkg::DISP_SIZE-1: 0] w_disp_grp_id;
  logic [msrh_pkg::LSU_INST_NUM-1: 0] w_ex2_ldq_entries_recv;

  for (genvar i_idx = 0; i_idx < msrh_conf_pkg::MEM_DISP_SIZE; i_idx++) begin : in_loop
    assign w_input_valid[i_idx] = disp_picked_inst_valid[i_idx] & (w_in_ptr + i_idx == l_idx);
  end

  bit_oh_or #(.WIDTH($size(msrh_pkg::disp_t)), .WORDS(msrh_conf_pkg::MEM_DISP_SIZE)) bit_oh_entry  (.i_oh(w_input_valid), .i_data(disp_picked_inst),   .o_selected(w_disp_entry));
  bit_oh_or #(.WIDTH(msrh_pkg::DISP_SIZE),     .WORDS(msrh_conf_pkg::MEM_DISP_SIZE)) bit_oh_grp_id (.i_oh(w_input_valid), .i_data(disp_picked_grp_id), .o_selected(w_disp_grp_id));

  // Selection of EX1 Update signal
  ex1_q_update_t w_ex1_q_updates;
  logic [msrh_pkg::LSU_INST_NUM-1: 0] w_ex1_q_valid;
  ex1_update_select u_ex1_update_select (.i_ex1_q_updates(i_ex1_q_updates), .cmt_id(w_ldq_entries[l_idx].cmt_id), .grp_id(w_ldq_entries[l_idx].grp_id),
                                         .o_ex1_q_valid(w_ex1_q_valid), .o_ex1_q_updates(w_ex1_q_updates));

  // Selection of EX1 Update signal
  ex2_q_update_t w_ex2_q_updates;
  logic w_ex2_q_valid;
  ex2_update_select u_ex2_update_select (.i_ex2_q_updates(i_ex2_q_updates),
                                         .q_index(l_idx[$clog2(LDQ_SIZE)-1:0]),
                                         .i_ex2_recv(w_ex2_ldq_entries_recv),
                                         .o_ex2_q_valid(w_ex2_q_valid), .o_ex2_q_updates(w_ex2_q_updates));

  msrh_ldq_entry
  u_msrh_ldq_entry
    (
     .i_clk     (i_clk    ),
     .i_reset_n (i_reset_n),

     .i_disp_load   (|w_input_valid),
     .i_disp_cmt_id (disp.cmt_id),
     .i_disp_grp_id (w_disp_grp_id),
     .i_disp        (w_disp_entry),

     .i_ex1_q_valid   (|w_ex1_q_valid),
     .i_ex1_q_updates (w_ex1_q_updates),

     .i_tlb_resolve (i_tlb_resolve),

     .i_ex2_q_valid  (|w_ex2_q_valid),
     .i_ex2_q_updates(w_ex2_q_updates),

     .o_entry (w_ldq_entries[l_idx]),
     .o_ex2_ldq_entries_recv(w_ex2_ldq_entries_recv),

     .i_rerun_accept (|w_rerun_request_rev_oh[l_idx] & !(|w_ldq_replay_conflict[l_idx])),

     .i_lrq_resolve (i_lrq_resolve),

     .i_ex3_done (i_ex3_done),
     .i_ldq_done (w_ldq_done_oh[l_idx])
     );

  for (genvar p_idx = 0; p_idx < msrh_pkg::LSU_INST_NUM; p_idx++) begin : pipe_loop
    assign w_rerun_request[p_idx][l_idx] = w_ldq_entries[l_idx].state == LDQ_READY &&
                                           w_ldq_entries[l_idx].pipe_sel_idx_oh[p_idx];
  end
end
endgenerate

// replay logic
generate for (genvar p_idx = 0; p_idx < msrh_pkg::LSU_INST_NUM; p_idx++) begin : pipe_loop
  assign ldq_replay_if[p_idx].valid = |w_rerun_request[p_idx];
  ldq_entry_t w_ldq_replay_entry;

  bit_extract_lsb #(.WIDTH(LDQ_SIZE)) u_bit_req_sel (.in(w_rerun_request[p_idx]), .out(w_rerun_request_oh[p_idx]));
  bit_oh_or #(.WIDTH($size(ldq_entry_t)), .WORDS(LDQ_SIZE)) select_rerun_oh  (.i_oh(w_rerun_request_oh[p_idx]), .i_data(w_ldq_entries), .o_selected(w_ldq_replay_entry));

  assign ldq_replay_if[p_idx].issue = w_ldq_replay_entry.inst;

  assign ldq_replay_if[p_idx].index_oh = w_rerun_request_oh[p_idx];

  for (genvar l_idx = 0; l_idx < LDQ_SIZE; l_idx++) begin : ldq_loop
    assign w_rerun_request_rev_oh[l_idx][p_idx] = w_rerun_request_oh[p_idx][l_idx];

    assign w_ldq_replay_conflict[l_idx][p_idx] = ldq_replay_if[p_idx].conflict & w_rerun_request[p_idx][l_idx];
  end
end
endgenerate

// ===============
// done logic
// ===============
generate for (genvar l_idx = 0; l_idx < LDQ_SIZE; l_idx++) begin : done_loop
  assign w_ldq_done_oh[l_idx] = w_ldq_entries[l_idx].state == LDQ_EX3_DONE && (w_out_ptr == l_idx);
end
endgenerate
bit_oh_or #(.WIDTH($size(ldq_entry_t)), .WORDS(LDQ_SIZE)) select_rerun_oh  (.i_oh(w_ldq_done_oh), .i_data(w_ldq_entries), .o_selected(w_ldq_done_entry));

assign o_done_report.valid   = |w_ldq_done_oh;
assign o_done_report.cmt_id  = w_ldq_done_entry.cmt_id;
assign o_done_report.grp_id  = w_ldq_done_entry.grp_id;
assign o_done_report.exc_vld = 'h0;   // Temporary

`ifdef SIMULATION

function void dump_entry_json(int fp, ldq_entry_t entry, int index);

  if (entry.is_valid) begin
    $fwrite(fp, "    \"msrh_ldq_entry[%d]\" : {", index);
    $fwrite(fp, "       valid : %d, ", entry.is_valid);
    $fwrite(fp, "       pc_addr : \"0x%0x\", ", entry.inst.pc_addr);
    $fwrite(fp, "       inst : \"%08x\", ", entry.inst);

    $fwrite(fp, "       cmt_id : %d, ", entry.cmt_id);
    $fwrite(fp, "       grp_id : %d, ", entry.grp_id);

    $fwrite(fp, "       state : \"%s\, ", entry.state == LDQ_INIT     ? "LDQ_INIT" :
                                          entry.state == LDQ_EX2_RUN  ? "LDQ_EX2_RUN" :
                                          entry.state == LDQ_LRQ_HAZ  ? "LDQ_LRQ_HAZ" :
                                          entry.state == LDQ_STQ_HAZ  ? "LDQ_STQ_HAZ" :
                                          entry.state == LDQ_TLB_HAZ  ? "LDQ_TLB_HAZ" :
                                          entry.state == LDQ_READY    ? "LDQ_READY" :
                                          entry.state == LDQ_EX3_DONE ? "LDQ_EX3_DONE" : "x");
    $fwrite(fp, "    },\n");
  end // if (entry.valid)

endfunction // dump_json

function void dump_json(int fp);
  $fwrite(fp, "  \"msrh_ldq\" : {\n");
  for (int l_idx = 0; l_idx < MEM_Q_SIZE; l_idx++) begin
    dump_entry_json (fp, w_ldq_entries[l_idx], l_idx);
  end
  $fwrite(fp, "  },\n");
endfunction // dump_json
`endif // SIMULATION

endmodule // msrh_ldq

module ex1_update_select
  import msrh_lsu_pkg::*;
  (
   input ex1_q_update_t i_ex1_q_updates[msrh_pkg::LSU_INST_NUM],
   input logic [msrh_pkg::CMT_BLK_W-1: 0] cmt_id,
   input logic [msrh_pkg::DISP_SIZE-1: 0] grp_id,
   output [msrh_pkg::LSU_INST_NUM-1: 0]   o_ex1_q_valid,
   output                                 ex1_q_update_t o_ex1_q_updates
   );

logic [msrh_pkg::LSU_INST_NUM-1: 0] w_ex1_update_match;

for (genvar p_idx = 0; p_idx < msrh_pkg::LSU_INST_NUM; p_idx++) begin : ex1_update_loop
  assign o_ex1_q_valid[p_idx] = i_ex1_q_updates[p_idx].update &&
                                i_ex1_q_updates[p_idx].cmt_id == cmt_id &&
                                i_ex1_q_updates[p_idx].grp_id == grp_id;
end

bit_oh_or #(.WIDTH($size(ex1_q_update_t)), .WORDS(msrh_pkg::LSU_INST_NUM)) bit_oh_update (.i_oh(o_ex1_q_valid), .i_data(i_ex1_q_updates), .o_selected(o_ex1_q_updates));

endmodule // ex1_update_select


module ex2_update_select
  import msrh_lsu_pkg::*;
  (
   input ex2_q_update_t i_ex2_q_updates[msrh_pkg::LSU_INST_NUM],
   input logic [$clog2(LDQ_SIZE)-1: 0] q_index,
   input logic [msrh_pkg::LSU_INST_NUM-1: 0]         i_ex2_recv,
   output                                            o_ex2_q_valid,
   output                                            ex2_q_update_t o_ex2_q_updates
   );

logic [msrh_pkg::LSU_INST_NUM-1: 0] w_ex2_update_match;

for (genvar p_idx = 0; p_idx < msrh_pkg::LSU_INST_NUM; p_idx++) begin : ex2_update_loop
  assign w_ex2_update_match[p_idx] = (i_ex2_q_updates[p_idx].update &&
                                      i_ex2_q_updates[p_idx].index_oh[q_index]) |
                                     i_ex2_recv[p_idx];
end

assign o_ex2_q_valid = |w_ex2_update_match;
bit_oh_or #(.WIDTH($size(ex2_q_update_t)), .WORDS(msrh_pkg::LSU_INST_NUM)) bit_oh_update (.i_oh(w_ex2_update_match), .i_data(i_ex2_q_updates), .o_selected(o_ex2_q_updates));

endmodule // ex2_update_select
