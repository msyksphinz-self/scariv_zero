riscv_fpu_imafdc_pkg.sv