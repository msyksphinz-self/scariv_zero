`define RV64
`define LITEX_SIMULATION
