// ------------------------------------------------------------------------
// NAME :
// TYPE : package
// ------------------------------------------------------------------------
//
// ------------------------------------------------------------------------
//
// ------------------------------------------------------------------------

interface br_upd_if;

  logic                                update;
  logic                                taken;
  logic                                mispredict;
  logic                                is_cond;
  logic                                is_call;
  logic                                is_ret;
  logic                                is_rvc;
  logic [$clog2(scariv_conf_pkg::RAS_ENTRY_SIZE)-1: 0] ras_index;
  logic [ 1: 0]                        bim_value;
  scariv_pkg::vaddr_t                    pc_vaddr;
  scariv_pkg::vaddr_t                    target_vaddr;
  scariv_pkg::vaddr_t                    ras_prev_vaddr;
`ifdef SIMULATION
  scariv_pkg::vaddr_t                    pred_vaddr;
`endif // SIMULATION
  logic                                dead;
  scariv_pkg::cmt_id_t                   cmt_id;
  scariv_pkg::grp_id_t                   grp_id;
  scariv_pkg::brtag_t                    brtag;

  logic [scariv_pkg::GSHARE_BHT_W-1: 0] gshare_index;
  logic [scariv_pkg::GSHARE_BHT_W-1: 0] gshare_bhr;

  modport master (
    output update,
    output taken,
    output mispredict,
    output is_cond,
    output is_call,
    output is_ret,
    output is_rvc,
    output ras_index,
    output bim_value,
    output dead,
    output pc_vaddr,
    output target_vaddr,
    output ras_prev_vaddr,
`ifdef SIMULATION
    output pred_vaddr,
`endif // SIMULATION
    output cmt_id,
    output grp_id,
    output brtag,
    output gshare_index,
    output gshare_bhr
  );

  modport slave (
    input update,
    input taken,
    input mispredict,
    input is_cond,
    input is_call,
    input is_ret,
    input is_rvc,
    input ras_index,
    input bim_value,
    input dead,
    input pc_vaddr,
    input target_vaddr,
    input ras_prev_vaddr,
`ifdef SIMULATION
    input pred_vaddr,
`endif // SIMULATION
    input cmt_id,
    input grp_id,
    input brtag,
    input gshare_index,
    input gshare_bhr
  );

endinterface // br_upd_if


module br_upd_if_buf
  (
   br_upd_if.slave  slave_if,
   br_upd_if.master master_if
   );

assign master_if.update         = slave_if.update         ;
assign master_if.taken          = slave_if.taken          ;
assign master_if.mispredict     = slave_if.mispredict     ;
assign master_if.is_cond        = slave_if.is_cond        ;
assign master_if.is_call        = slave_if.is_call        ;
assign master_if.is_ret         = slave_if.is_ret         ;
assign master_if.is_rvc         = slave_if.is_rvc         ;
assign master_if.ras_index      = slave_if.ras_index      ;
assign master_if.bim_value      = slave_if.bim_value      ;
assign master_if.pc_vaddr       = slave_if.pc_vaddr       ;
assign master_if.target_vaddr   = slave_if.target_vaddr   ;
assign master_if.ras_prev_vaddr = slave_if.ras_prev_vaddr ;
`ifdef SIMULATION
assign master_if.pred_vaddr     = slave_if.pred_vaddr     ;
`endif // SIMULATION
assign master_if.dead           = slave_if.dead           ;
assign master_if.cmt_id         = slave_if.cmt_id         ;
assign master_if.grp_id         = slave_if.grp_id         ;
assign master_if.brtag          = slave_if.brtag          ;
assign master_if.gshare_index   = slave_if.gshare_index    ;
assign master_if.gshare_bhr     = slave_if.gshare_bhr      ;

endmodule // br_upd_if_buf


interface cmt_brtag_if;

  logic          commit;
  scariv_pkg::grp_id_t is_br_inst;
  logic [scariv_conf_pkg::DISP_SIZE-1: 0][$clog2(scariv_conf_pkg::RV_BRU_ENTRY_SIZE)-1: 0] brtag;
  scariv_pkg::gshare_bht_t gshare_bhr;
  scariv_pkg::gshare_bht_t gshare_index;
  logic                    taken;
  logic [ 1: 0]            bim_value;
  logic                    is_rvc;
  logic                    dead;

  modport master (
    output commit,
    output is_br_inst,
    output brtag,
    output gshare_bhr,
    output gshare_index,
    output taken,
    output bim_value,
    output is_rvc,
    output dead
  );

  modport slave (
    input commit,
    input is_br_inst,
    input brtag,
    input gshare_bhr,
    input gshare_index,
    input taken,
    input bim_value,
    input is_rvc,
    input dead
  );

endinterface // cmt_brtag_if

interface brtag_if;
  logic valid;
  scariv_pkg::brtag_t brtag;

  modport master (
    output valid,
    output brtag
  );

  modport slave (
    input valid,
    input brtag
  );
endinterface
