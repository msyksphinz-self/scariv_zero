// ------------------------------------------------------------------------
// NAME : scariv_fpu_pkg
// TYPE : package
// ------------------------------------------------------------------------
// FPU Package
// ------------------------------------------------------------------------
// ------------------------------------------------------------------------

package scariv_fpu_pkg;

import decoder_fpu_ctrl_pkg::*;

endpackage // scariv_fpu_pkg
