`default_nettype none

package riscv_pkg;

  localparam XLEN_W = 64;
  localparam PADDR_W = 39;

endpackage

`default_nettype wire
