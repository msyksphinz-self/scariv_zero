// Generator : SpinalHDL dev    git head : 700e223f5dc8c2258117fae140ab8d6eb8446d97
// Component : NaxRiscv
// Git hash  : 3fa251104e4bc3cb5fda8e784838fd94200875d6

`timescale 1ns/1ps

module NaxRiscv (
  output wire          FetchCachePlugin_mem_cmd_valid,
  input  wire          FetchCachePlugin_mem_cmd_ready,
  output wire [31:0]   FetchCachePlugin_mem_cmd_payload_address,
  output wire          FetchCachePlugin_mem_cmd_payload_io,
  input  wire          FetchCachePlugin_mem_rsp_valid,
  output wire          FetchCachePlugin_mem_rsp_ready,
  input  wire [63:0]   FetchCachePlugin_mem_rsp_payload_data,
  input  wire          FetchCachePlugin_mem_rsp_payload_error,
  input  wire          PrivilegedPlugin_io_int_machine_timer /* verilator public */ ,
  input  wire          PrivilegedPlugin_io_int_machine_software /* verilator public */ ,
  input  wire          PrivilegedPlugin_io_int_machine_external /* verilator public */ ,
  input  wire          PrivilegedPlugin_io_int_supervisor_external /* verilator public */ ,
  input  wire [63:0]   PrivilegedPlugin_io_rdtime,
  output wire          LsuPlugin_peripheralBus_cmd_valid /* verilator public */ ,
  input  wire          LsuPlugin_peripheralBus_cmd_ready /* verilator public */ ,
  output wire          LsuPlugin_peripheralBus_cmd_payload_write /* verilator public */ ,
  output wire [31:0]   LsuPlugin_peripheralBus_cmd_payload_address /* verilator public */ ,
  output wire [31:0]   LsuPlugin_peripheralBus_cmd_payload_data /* verilator public */ ,
  output wire [3:0]    LsuPlugin_peripheralBus_cmd_payload_mask /* verilator public */ ,
  output wire [1:0]    LsuPlugin_peripheralBus_cmd_payload_size /* verilator public */ ,
  input  wire          LsuPlugin_peripheralBus_rsp_valid /* verilator public */ ,
  input  wire          LsuPlugin_peripheralBus_rsp_payload_error /* verilator public */ ,
  input  wire [31:0]   LsuPlugin_peripheralBus_rsp_payload_data /* verilator public */ ,
  output wire          DataCachePlugin_mem_read_cmd_valid,
  input  wire          DataCachePlugin_mem_read_cmd_ready,
  output wire [0:0]    DataCachePlugin_mem_read_cmd_payload_id,
  output wire [31:0]   DataCachePlugin_mem_read_cmd_payload_address,
  input  wire          DataCachePlugin_mem_read_rsp_valid,
  output wire          DataCachePlugin_mem_read_rsp_ready,
  input  wire [0:0]    DataCachePlugin_mem_read_rsp_payload_id,
  input  wire [63:0]   DataCachePlugin_mem_read_rsp_payload_data,
  input  wire          DataCachePlugin_mem_read_rsp_payload_error,
  output wire          DataCachePlugin_mem_write_cmd_valid,
  input  wire          DataCachePlugin_mem_write_cmd_ready,
  output wire          DataCachePlugin_mem_write_cmd_payload_last,
  output wire [31:0]   DataCachePlugin_mem_write_cmd_payload_fragment_address,
  output wire [63:0]   DataCachePlugin_mem_write_cmd_payload_fragment_data,
  output wire [0:0]    DataCachePlugin_mem_write_cmd_payload_fragment_id,
  input  wire          DataCachePlugin_mem_write_rsp_valid,
  input  wire          DataCachePlugin_mem_write_rsp_payload_error,
  input  wire [0:0]    DataCachePlugin_mem_write_rsp_payload_id,
  input  wire          clk,
  input  wire          reset
);
  localparam BranchPlugin_BranchCtrlEnum_B = 2'd0;
  localparam BranchPlugin_BranchCtrlEnum_JAL = 2'd1;
  localparam BranchPlugin_BranchCtrlEnum_JALR = 2'd2;
  localparam IntAluPlugin_AluCtrlEnum_ADD_SUB = 2'd0;
  localparam IntAluPlugin_AluCtrlEnum_SLT_SLTU = 2'd1;
  localparam IntAluPlugin_AluCtrlEnum_BITWISE = 2'd2;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 = 2'd0;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_OR_1 = 2'd1;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_AND_1 = 2'd2;
  localparam Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN = 3'd0;
  localparam Lsu2Plugin_CTRL_ENUM_MMU_REDO = 3'd1;
  localparam Lsu2Plugin_CTRL_ENUM_TRAP_MMU = 3'd2;
  localparam Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD = 3'd3;
  localparam Lsu2Plugin_CTRL_ENUM_LOAD_MISS = 3'd4;
  localparam Lsu2Plugin_CTRL_ENUM_LOAD_FAILED = 3'd5;
  localparam Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS = 3'd6;
  localparam Lsu2Plugin_CTRL_ENUM_SUCCESS = 3'd7;
  localparam EnvCallPlugin_logic_flushes_enumDef_BOOT = 3'd0;
  localparam EnvCallPlugin_logic_flushes_enumDef_IDLE = 3'd1;
  localparam EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE = 3'd2;
  localparam EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH = 3'd3;
  localparam EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT = 3'd4;
  localparam EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH = 3'd5;
  localparam EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU = 3'd6;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_BOOT = 9'd1;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_IDLE = 9'd2;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD = 9'd4;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP = 9'd8;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY = 9'd16;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_ALU = 9'd32;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION = 9'd64;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_SYNC = 9'd128;
  localparam Lsu2Plugin_logic_special_atomic_enumDef_TRAP = 9'd256;
  localparam PrivilegedPlugin_logic_fsm_enumDef_BOOT = 4'd0;
  localparam PrivilegedPlugin_logic_fsm_enumDef_IDLE = 4'd1;
  localparam PrivilegedPlugin_logic_fsm_enumDef_SETUP = 4'd2;
  localparam PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE = 4'd3;
  localparam PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE = 4'd4;
  localparam PrivilegedPlugin_logic_fsm_enumDef_EPC_READ = 4'd5;
  localparam PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ = 4'd6;
  localparam PrivilegedPlugin_logic_fsm_enumDef_XRET = 4'd7;
  localparam PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC = 4'd8;
  localparam PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP = 4'd9;
  localparam PrivilegedPlugin_logic_fsm_enumDef_TRAP = 4'd10;
  localparam MmuPlugin_logic_refill_enumDef_BOOT = 3'd0;
  localparam MmuPlugin_logic_refill_enumDef_IDLE = 3'd1;
  localparam MmuPlugin_logic_refill_enumDef_INIT = 3'd2;
  localparam MmuPlugin_logic_refill_enumDef_CMD_0 = 3'd3;
  localparam MmuPlugin_logic_refill_enumDef_CMD_1 = 3'd4;
  localparam MmuPlugin_logic_refill_enumDef_RSP_0 = 3'd5;
  localparam MmuPlugin_logic_refill_enumDef_RSP_1 = 3'd6;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT = 3'd0;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE = 3'd1;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_READ = 3'd2;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE = 3'd3;
  localparam EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE = 3'd4;
  localparam PerformanceCounterPlugin_logic_fsm_enumDef_BOOT = 4'd0;
  localparam PerformanceCounterPlugin_logic_fsm_enumDef_IDLE = 4'd1;
  localparam PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW = 4'd2;
  localparam PerformanceCounterPlugin_logic_fsm_enumDef_CALC = 4'd3;
  localparam PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW = 4'd4;
  localparam PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH = 4'd5;
  localparam PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH = 4'd6;
  localparam PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE = 4'd7;
  localparam PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION = 4'd8;

  reg                 integer_RfTranslationPlugin_logic_impl_io_rollback;
  wire                integer_RfTranslationPlugin_logic_impl_io_writes_0_valid;
  wire                integer_RfTranslationPlugin_logic_impl_io_writes_1_valid;
  reg                 integer_RfTranslationPlugin_logic_impl_io_commits_0_valid;
  reg        [4:0]    integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_address;
  reg        [5:0]    integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_data;
  wire                integer_RfTranslationPlugin_logic_impl_io_commits_1_valid;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_0_cmd_valid;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_1_cmd_valid;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_2_cmd_valid;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_3_cmd_valid;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_4_cmd_valid;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_5_cmd_valid;
  reg                 integer_RfAllocationPlugin_logic_allocator_io_push_0_valid;
  reg        [5:0]    integer_RfAllocationPlugin_logic_allocator_io_push_0_payload;
  reg                 integer_RfAllocationPlugin_logic_allocator_io_push_1_valid;
  wire       [5:0]    integer_RfAllocationPlugin_logic_allocator_io_push_1_payload;
  reg        [1:0]    integer_RfAllocationPlugin_logic_allocator_io_pop_mask;
  wire       [31:0]   DataCachePlugin_logic_cache_io_load_cmd_payload_virtual;
  wire       [1:0]    DataCachePlugin_logic_cache_io_load_cmd_payload_size;
  wire                DataCachePlugin_logic_cache_io_load_cmd_payload_redoOnDataHazard;
  wire                DataCachePlugin_logic_cache_io_load_cmd_payload_unlocked;
  wire                DataCachePlugin_logic_cache_io_load_cmd_payload_unique;
  wire       [31:0]   DataCachePlugin_logic_cache_io_load_translated_physical;
  wire                DataCachePlugin_logic_cache_io_load_translated_abord;
  wire       [2:0]    DataCachePlugin_logic_cache_io_load_cancels;
  wire                CommitPlugin_logic_free_lineEventStream_fifo_io_pop_ready;
  wire                CommitPlugin_logic_free_lineEventStream_fifo_io_flush;
  wire                EU0_DivPlugin_logic_div_io_cmd_valid;
  reg                 Lsu2Plugin_logic_prefetch_predictor_io_learn_valid;
  reg                 Lsu2Plugin_logic_prefetch_predictor_io_learn_payload_allocate;
  reg                 Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready;
  wire                Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_valid;
  wire                Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_payload;
  wire       [31:0]   DispatchPlugin_logic_queue_io_push_payload_slots_0_event;
  wire       [1:0]    DispatchPlugin_logic_queue_io_push_payload_slots_0_sel;
  wire       [0:0]    DispatchPlugin_logic_queue_io_push_payload_slots_0_context_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_push_payload_slots_0_context_robId;
  wire       [31:0]   DispatchPlugin_logic_queue_io_push_payload_slots_1_event;
  wire       [1:0]    DispatchPlugin_logic_queue_io_push_payload_slots_1_sel;
  wire       [0:0]    DispatchPlugin_logic_queue_io_push_payload_slots_1_context_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_push_payload_slots_1_context_robId;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_valid;
  wire       [5:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_payload_robId;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_writes_1_valid;
  wire       [5:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_writes_1_payload_robId;
  reg                 RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_valid;
  reg        [5:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_payload_physical;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_commits_1_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_commits_2_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_commits_3_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_commits_4_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_commits_5_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_cmd_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_cmd_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_cmd_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_cmd_valid;
  wire       [32:0]   BranchContextPlugin_logic_mem_earlyBranch_io_writes_0_payload_data;
  wire       [32:0]   BranchContextPlugin_logic_mem_earlyBranch_io_writes_1_payload_data;
  wire                BranchContextPlugin_logic_mem_earlyBranch_io_read_0_cmd_valid;
  wire                BranchContextPlugin_logic_mem_earlyBranch_io_read_1_cmd_valid;
  wire       [64:0]   BranchContextPlugin_logic_mem_finalBranch_io_writes_0_payload_data;
  wire       [64:0]   BranchContextPlugin_logic_mem_finalBranch_io_writes_1_payload_data;
  wire                BranchContextPlugin_logic_mem_finalBranch_io_read_0_cmd_valid;
  wire       [4:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_io_writes_0_payload_data;
  wire       [4:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_io_writes_1_payload_data;
  wire                Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_0_cmd_valid;
  wire                Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_1_cmd_valid;
  wire       [3:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_1_cmd_payload;
  wire                Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_2_cmd_valid;
  wire                Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_3_cmd_valid;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_doSpecial_io_writes_0_payload_data;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_doSpecial_io_writes_1_payload_data;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_doSpecial_io_writes_2_payload_data;
  wire                Lsu2Plugin_logic_lq_mem_doSpecial_io_read_0_cmd_valid;
  wire       [3:0]    Lsu2Plugin_logic_lq_mem_needTranslation_io_writes_0_payload_address;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_needTranslation_io_writes_0_payload_data;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_needTranslation_io_writes_1_payload_data;
  wire                Lsu2Plugin_logic_lq_mem_needTranslation_io_read_0_cmd_valid;
  wire       [3:0]    Lsu2Plugin_logic_sq_mem_needTranslation_io_writes_0_payload_address;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_needTranslation_io_writes_0_payload_data;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_needTranslation_io_writes_1_payload_data;
  wire                Lsu2Plugin_logic_sq_mem_needTranslation_io_read_0_cmd_valid;
  wire                Lsu2Plugin_logic_sq_mem_needTranslation_io_read_1_cmd_valid;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_feededOnce_io_writes_0_payload_data;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_feededOnce_io_writes_1_payload_data;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_feededOnce_io_writes_2_payload_data;
  wire                Lsu2Plugin_logic_sq_mem_feededOnce_io_read_0_cmd_valid;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_doSpecial_io_writes_0_payload_data;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_doSpecial_io_writes_1_payload_data;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_doSpecial_io_writes_2_payload_data;
  wire                Lsu2Plugin_logic_sq_mem_doSpecial_io_read_0_cmd_valid;
  wire       [4:0]    Lsu2Plugin_logic_sq_mem_lqAlloc_io_writes_0_payload_data;
  wire       [4:0]    Lsu2Plugin_logic_sq_mem_lqAlloc_io_writes_1_payload_data;
  wire                Lsu2Plugin_logic_sq_mem_lqAlloc_io_read_0_cmd_valid;
  wire                BranchContextPlugin_free_dispatchMem_mem_io_read_0_cmd_valid;
  wire                RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_0_valid;
  wire       [0:0]    RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_0_payload_data;
  wire                RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_1_valid;
  wire       [0:0]    RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_1_payload_data;
  wire                RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_0_cmd_valid;
  wire       [5:0]    RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_0_cmd_payload;
  wire                RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_1_cmd_valid;
  wire       [5:0]    RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_1_cmd_payload;
  wire                RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_2_cmd_valid;
  reg        [63:0]   _zz_FetchCachePlugin_logic_banks_0_mem_port1;
  reg        [63:0]   _zz_FetchCachePlugin_logic_banks_1_mem_port1;
  reg        [63:0]   _zz_FetchCachePlugin_logic_banks_2_mem_port1;
  reg        [63:0]   _zz_FetchCachePlugin_logic_banks_3_mem_port1;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_0_mem_port1;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_1_mem_port1;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_2_mem_port1;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_3_mem_port1;
  wire       [2:0]    _zz_FetchCachePlugin_logic_plru_ram_port1;
  wire       [31:0]   _zz_DecoderPredictionPlugin_logic_ras_mem_stack_port0;
  reg        [49:0]   _zz_BtbPlugin_logic_mem_port1;
  reg        [3:0]    _zz_GSharePlugin_logic_mem_counter_port1;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_addressPre_port1;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_addressPre_port2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_addressPost_port0;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_addressPost_port2;
  wire       [1:0]    _zz_Lsu2Plugin_logic_lq_mem_size_port1;
  wire       [1:0]    _zz_Lsu2Plugin_logic_lq_mem_size_port2;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_physRd_port1;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_physRd_port2;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_robId_port1;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_robId_port2;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_robId_port3;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port1;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_pc_port1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_io_port0;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_writeRd_port1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_writeRd_port2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_lr_port1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_unsigned_port1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_unsigned_port2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port1;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port1;
  reg        [22:0]   _zz_Lsu2Plugin_logic_lq_hazardPrediction_mem_port1;
  reg        [5:0]    _zz_Lsu2Plugin_logic_lq_hitPrediction_mem_port1;
  wire       [5:0]    _zz_Lsu2Plugin_logic_sq_mem_robId_port1;
  wire       [5:0]    _zz_Lsu2Plugin_logic_sq_mem_robId_port2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port1;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_addressPre_port1;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_addressPre_port2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_addressPost_port0;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_addressPost_port2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_addressPost_port3;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sq_mem_size_port1;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sq_mem_size_port2;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sq_mem_size_port3;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sq_mem_size_port4;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_io_port0;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_io_port2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_amo_port1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_amo_port2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_sc_port1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_sc_port2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_data_port1;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_data_port2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port1;
  wire       [41:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port1;
  wire       [41:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port1;
  wire       [41:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port1;
  wire       [41:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port1;
  wire       [21:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port1;
  wire       [21:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port1;
  wire       [41:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port1;
  wire       [41:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port1;
  wire       [41:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port1;
  wire       [41:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port1;
  wire       [21:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port1;
  wire       [21:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port1;
  wire       [31:0]   _zz_CsrRamPlugin_logic_mem_port1;
  wire       [1:0]    _zz_RobPlugin_logic_completionMem_target_port1;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_0_port0;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_0_port1;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_0_port2;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_0_port4;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_0_port5;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_1_port0;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_1_port1;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_1_port2;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_1_port4;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_1_port5;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_2_port0;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_2_port1;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_2_port2;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_2_port4;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_2_port5;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_3_port0;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_3_port1;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_3_port2;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_3_port4;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_3_port5;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_4_port0;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_4_port1;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_4_port2;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_4_port4;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_4_port5;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_5_port0;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_5_port1;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_5_port2;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_5_port4;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_5_port5;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_6_port0;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_6_port1;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_6_port2;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_6_port4;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_6_port5;
  wire       [1:0]    _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port1;
  wire       [1:0]    _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port2;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_0_port1;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_0_port2;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_0_port3;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_0_port4;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_1_port1;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_1_port2;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_1_port3;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_1_port4;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port3;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port4;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port3;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port4;
  wire       [11:0]   _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port1;
  wire       [11:0]   _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port2;
  wire       [9:0]    _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port1;
  wire       [11:0]   _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port1;
  wire       [1:0]    _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port2;
  wire       [23:0]   _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_port1;
  wire       [23:0]   _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_1_port1;
  wire       [3:0]    _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port1;
  wire       [3:0]    _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1_port1;
  wire       [1:0]    _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port1;
  wire       [1:0]    _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port1;
  wire       [31:0]   _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port1;
  wire       [31:0]   _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port2;
  wire       [31:0]   _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1_port1;
  wire       [31:0]   _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1_port2;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port1;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_1_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port2;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port1;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_1_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port2;
  wire       [3:0]    _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port1;
  wire       [3:0]    _zz_RobPlugin_logic_storage_BRANCH_ID_banks_1_port1;
  wire       [4:0]    _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port1;
  wire       [4:0]    _zz_RobPlugin_logic_storage_LSU_ID_banks_1_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_ROB_MSB_banks_1_port1;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_valid;
  wire       [5:0]    integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_payload;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_valid;
  wire       [5:0]    integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_payload;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_valid;
  wire       [5:0]    integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_payload;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_3_rsp_valid;
  wire       [5:0]    integer_RfTranslationPlugin_logic_impl_io_reads_3_rsp_payload;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_4_rsp_valid;
  wire       [5:0]    integer_RfTranslationPlugin_logic_impl_io_reads_4_rsp_payload;
  wire                integer_RfTranslationPlugin_logic_impl_io_reads_5_rsp_valid;
  wire       [5:0]    integer_RfTranslationPlugin_logic_impl_io_reads_5_rsp_payload;
  wire                integer_RfAllocationPlugin_logic_allocator_io_pop_ready;
  wire       [5:0]    integer_RfAllocationPlugin_logic_allocator_io_pop_values_0;
  wire       [5:0]    integer_RfAllocationPlugin_logic_allocator_io_pop_values_1;
  wire                DataCachePlugin_logic_cache_io_load_cmd_ready;
  wire                DataCachePlugin_logic_cache_io_load_rsp_valid;
  wire       [31:0]   DataCachePlugin_logic_cache_io_load_rsp_payload_data;
  wire                DataCachePlugin_logic_cache_io_load_rsp_payload_fault;
  wire                DataCachePlugin_logic_cache_io_load_rsp_payload_redo;
  wire       [1:0]    DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlot;
  wire                DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlotAny;
  wire                DataCachePlugin_logic_cache_io_store_cmd_ready;
  wire                DataCachePlugin_logic_cache_io_store_rsp_valid;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_fault;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_redo;
  wire       [1:0]    DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlot;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlotAny;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_generationKo;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_flush;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_prefetch;
  wire       [31:0]   DataCachePlugin_logic_cache_io_store_rsp_payload_address;
  wire                DataCachePlugin_logic_cache_io_store_rsp_payload_io;
  wire                DataCachePlugin_logic_cache_io_mem_read_cmd_valid;
  wire       [0:0]    DataCachePlugin_logic_cache_io_mem_read_cmd_payload_id;
  wire       [31:0]   DataCachePlugin_logic_cache_io_mem_read_cmd_payload_address;
  wire                DataCachePlugin_logic_cache_io_mem_read_rsp_ready;
  wire                DataCachePlugin_logic_cache_io_mem_write_cmd_valid;
  wire                DataCachePlugin_logic_cache_io_mem_write_cmd_payload_last;
  wire       [31:0]   DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_address;
  wire       [63:0]   DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_data;
  wire       [0:0]    DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_id;
  wire       [1:0]    DataCachePlugin_logic_cache_io_refillCompletions;
  wire                DataCachePlugin_logic_cache_io_refillEvent;
  wire                DataCachePlugin_logic_cache_io_writebackEvent;
  wire                DataCachePlugin_logic_cache_io_writebackBusy;
  wire                DataCachePlugin_logic_cache_io_tagEvent;
  wire                CommitPlugin_logic_free_lineEventStream_fifo_io_push_ready;
  wire                CommitPlugin_logic_free_lineEventStream_fifo_io_pop_valid;
  wire       [5:0]    CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_robId;
  wire       [1:0]    CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_mask;
  wire       [5:0]    CommitPlugin_logic_free_lineEventStream_fifo_io_occupancy;
  wire       [5:0]    CommitPlugin_logic_free_lineEventStream_fifo_io_availability;
  wire                EU0_DivPlugin_logic_div_io_cmd_ready;
  wire                EU0_DivPlugin_logic_div_io_rsp_valid;
  wire       [34:0]   EU0_DivPlugin_logic_div_io_rsp_payload_result;
  wire       [32:0]   EU0_DivPlugin_logic_div_io_rsp_payload_remain;
  wire                Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_valid;
  wire       [31:0]   Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_payload;
  wire                DispatchPlugin_logic_queue_io_push_ready;
  wire                DispatchPlugin_logic_queue_io_schedules_0_valid;
  wire       [15:0]   DispatchPlugin_logic_queue_io_schedules_0_payload_event;
  wire                DispatchPlugin_logic_queue_io_schedules_1_valid;
  wire       [15:0]   DispatchPlugin_logic_queue_io_schedules_1_payload_event;
  wire                DispatchPlugin_logic_queue_io_schedules_2_valid;
  wire       [31:0]   DispatchPlugin_logic_queue_io_schedules_2_payload_event;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_0_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_0_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_0_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_0_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_0_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_1_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_1_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_1_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_1_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_1_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_2_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_2_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_2_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_2_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_2_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_3_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_3_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_3_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_3_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_3_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_4_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_4_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_4_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_4_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_4_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_5_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_5_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_5_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_5_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_5_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_6_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_6_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_6_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_6_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_6_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_7_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_7_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_7_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_7_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_7_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_8_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_8_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_8_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_8_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_8_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_9_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_9_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_9_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_9_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_9_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_10_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_10_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_10_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_10_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_10_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_11_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_11_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_11_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_11_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_11_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_12_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_12_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_12_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_12_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_12_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_13_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_13_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_13_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_13_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_13_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_14_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_14_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_14_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_14_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_14_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_15_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_15_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_15_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_15_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_15_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_16_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_16_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_16_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_16_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_16_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_17_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_17_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_17_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_17_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_17_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_18_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_18_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_18_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_18_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_18_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_19_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_19_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_19_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_19_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_19_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_20_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_20_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_20_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_20_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_20_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_21_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_21_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_21_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_21_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_21_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_22_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_22_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_22_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_22_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_22_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_23_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_23_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_23_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_23_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_23_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_24_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_24_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_24_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_24_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_24_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_25_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_25_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_25_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_25_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_25_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_26_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_26_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_26_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_26_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_26_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_27_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_27_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_27_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_27_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_27_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_28_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_28_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_28_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_28_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_28_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_29_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_29_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_29_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_29_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_29_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_30_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_30_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_30_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_30_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_30_euCtx_1;
  wire       [0:0]    DispatchPlugin_logic_queue_io_contexts_31_staticWake;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_31_physRd;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_31_robId;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_31_euCtx_0;
  wire       [5:0]    DispatchPlugin_logic_queue_io_contexts_31_euCtx_1;
  wire       [31:0]   DispatchPlugin_logic_queue_io_usage;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_2_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_3_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_4_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_5_data;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_enable;
  wire       [5:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_rob;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_enable;
  wire       [5:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_rob;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_rsp_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_rsp_payload_enable;
  wire       [5:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_rsp_payload_rob;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_rsp_valid;
  wire                RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_rsp_payload_enable;
  wire       [5:0]    RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_rsp_payload_rob;
  wire       [32:0]   BranchContextPlugin_logic_mem_earlyBranch_io_read_0_rsp;
  wire       [32:0]   BranchContextPlugin_logic_mem_earlyBranch_io_read_1_rsp;
  wire       [64:0]   BranchContextPlugin_logic_mem_finalBranch_io_read_0_rsp;
  wire       [4:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_0_rsp;
  wire       [4:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_1_rsp;
  wire       [4:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_2_rsp;
  wire       [4:0]    Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_3_rsp;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_doSpecial_io_read_0_rsp;
  wire       [0:0]    Lsu2Plugin_logic_lq_mem_needTranslation_io_read_0_rsp;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_needTranslation_io_read_0_rsp;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_needTranslation_io_read_1_rsp;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_feededOnce_io_read_0_rsp;
  wire       [0:0]    Lsu2Plugin_logic_sq_mem_doSpecial_io_read_0_rsp;
  wire       [4:0]    Lsu2Plugin_logic_sq_mem_lqAlloc_io_read_0_rsp;
  wire       [28:0]   BranchContextPlugin_free_dispatchMem_mem_io_read_0_rsp;
  wire       [0:0]    RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_0_rsp;
  wire       [0:0]    RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_1_rsp;
  wire       [0:0]    RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_2_rsp;
  wire       [11:0]   _zz_FetchPlugin_stages_1_FETCH_ID;
  wire       [0:0]    _zz_FetchPlugin_stages_1_FETCH_ID_1;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_0_mem_port;
  wire                _zz_FetchCachePlugin_logic_ways_0_mem_port_1;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_1_mem_port;
  wire                _zz_FetchCachePlugin_logic_ways_1_mem_port_1;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_2_mem_port;
  wire                _zz_FetchCachePlugin_logic_ways_2_mem_port_1;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_3_mem_port;
  wire                _zz_FetchCachePlugin_logic_ways_3_mem_port_1;
  wire       [2:0]    _zz_FetchCachePlugin_logic_plru_ram_port;
  wire       [1:0]    _zz_FetchCachePlugin_logic_refill_randomWay_valueNext;
  wire       [0:0]    _zz_FetchCachePlugin_logic_refill_randomWay_valueNext_1;
  wire       [19:0]   _zz_FetchCachePlugin_logic_read_onWays_0_hits_bypassHits;
  wire       [19:0]   _zz_FetchCachePlugin_logic_read_onWays_1_hits_bypassHits;
  wire       [19:0]   _zz_FetchCachePlugin_logic_read_onWays_2_hits_bypassHits;
  wire       [19:0]   _zz_FetchCachePlugin_logic_read_onWays_3_hits_bypassHits;
  reg        [1:0]    _zz_FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT;
  wire       [0:0]    _zz_FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT_1;
  reg        [1:0]    _zz_AlignerPlugin_setup_s2m_MASK_BACK;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_usable;
  reg        [31:0]   _zz_AlignerPlugin_logic_extractors_0_pcWord;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_pcWord_1;
  wire       [28:0]   _zz_FrontendPlugin_aligned_PC_0;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_usable;
  reg        [31:0]   _zz_AlignerPlugin_logic_extractors_1_pcWord;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_1_pcWord_1;
  wire       [28:0]   _zz_FrontendPlugin_aligned_PC_1;
  wire       [1:0]    _zz_DispatchPlugin_logic_sparseRob_sparse_ohFirst_masked;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push_1;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push_2;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push_3;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_push_4;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_1;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_2;
  wire       [3:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_3;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_4;
  wire       [31:0]   _zz_DecoderPredictionPlugin_logic_ras_mem_stack_port;
  wire       [49:0]   _zz_BtbPlugin_logic_mem_port;
  wire       [28:0]   _zz_BtbPlugin_logic_onLearn_port_payload_address;
  wire       [29:0]   _zz_BtbPlugin_logic_onLearn_port_payload_data_slice;
  wire       [28:0]   _zz_BtbPlugin_logic_readCmd_entryAddress;
  reg                 _zz_BtbPlugin_logic_applyIt_prediction;
  wire       [3:0]    _zz_GSharePlugin_logic_mem_counter_port;
  wire                _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_1;
  wire       [0:0]    _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_2;
  wire       [4:0]    _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_3;
  wire       [12:0]   _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_4;
  wire       [23:0]   _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_5;
  wire                _zz_GSharePlugin_logic_onLearn_hash_1;
  wire       [0:0]    _zz_GSharePlugin_logic_onLearn_hash_2;
  wire       [4:0]    _zz_GSharePlugin_logic_onLearn_hash_3;
  wire       [12:0]   _zz_GSharePlugin_logic_onLearn_hash_4;
  wire       [23:0]   _zz_GSharePlugin_logic_onLearn_hash_5;
  wire       [6:0]    _zz_CommitPlugin_logic_ptr_allocNext;
  wire       [1:0]    _zz_CommitPlugin_logic_ptr_allocNext_1;
  wire       [4:0]    _zz_CommitPlugin_logic_reschedule_commit_rowHit;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_age;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_0_age;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_1_age;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_2_age;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_3_age;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_4_age;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_5_age;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_1;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_2;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_3;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_4;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_5;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_6;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_7;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_8;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_9;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_10;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_11;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_12;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_13;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_14;
  wire                _zz_CommitPlugin_logic_reschedule_portsLogic_hits_15;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_robId;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_robId_1;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_robId_2;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_robId_3;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_robId_4;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_robId_5;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_robId_6;
  wire       [5:0]    _zz_CommitPlugin_logic_reschedule_robId_7;
  wire       [0:0]    _zz_CommitPlugin_logic_reschedule_trap_6;
  wire                _zz_CommitPlugin_logic_reschedule_cause;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_cause_1;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_cause_2;
  wire                _zz_CommitPlugin_logic_reschedule_cause_3;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_cause_4;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_cause_5;
  wire                _zz_CommitPlugin_logic_reschedule_cause_6;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_cause_7;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_cause_8;
  wire                _zz_CommitPlugin_logic_reschedule_cause_9;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_cause_10;
  wire       [3:0]    _zz_CommitPlugin_logic_reschedule_cause_11;
  wire                _zz_CommitPlugin_logic_reschedule_reason;
  wire       [7:0]    _zz_CommitPlugin_logic_reschedule_reason_1;
  wire       [7:0]    _zz_CommitPlugin_logic_reschedule_reason_2;
  wire                _zz_CommitPlugin_logic_reschedule_reason_3;
  wire       [7:0]    _zz_CommitPlugin_logic_reschedule_reason_4;
  wire       [7:0]    _zz_CommitPlugin_logic_reschedule_reason_5;
  wire                _zz_CommitPlugin_logic_reschedule_reason_6;
  wire       [7:0]    _zz_CommitPlugin_logic_reschedule_reason_7;
  wire       [7:0]    _zz_CommitPlugin_logic_reschedule_reason_8;
  wire                _zz_CommitPlugin_logic_reschedule_reason_9;
  wire       [7:0]    _zz_CommitPlugin_logic_reschedule_reason_10;
  wire       [7:0]    _zz_CommitPlugin_logic_reschedule_reason_11;
  wire       [0:0]    _zz_CommitPlugin_logic_reschedule_skipCommit;
  wire       [1:0]    _zz__zz_CommitPlugin_logic_commit_head_1;
  wire       [1:0]    _zz__zz_CommitPlugin_logic_commit_head_1_1;
  wire       [6:0]    _zz_CommitPlugin_logic_commit_head_2;
  wire       [6:0]    _zz_CommitPlugin_logic_commit_head_3;
  wire       [0:0]    _zz_CommitPlugin_logic_commit_head_4;
  wire       [5:0]    _zz_CommitPlugin_logic_free_robHit;
  reg        [1:0]    _zz_CommitDebugFilterPlugin_logic_commits_2;
  wire       [1:0]    _zz_CommitDebugFilterPlugin_logic_commits_3;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_0_value;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_0_value_1;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_0_value_2;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_0_value_3;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_1_value;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_1_value_1;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_1_value_2;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_1_value_3;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_2_value;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_2_value_1;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_2_value_2;
  wire       [31:0]   _zz_CommitDebugFilterPlugin_logic_filters_2_value_3;
  reg        [31:0]   _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_2;
  wire       [0:0]    _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_3;
  reg        [1:0]    _zz_PerformanceCounterPlugin_logic_commitCount;
  wire       [1:0]    _zz_PerformanceCounterPlugin_logic_commitCount_1;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_0;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_0_1;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_1_1;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_2;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_2_1;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_3;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_3_1;
  wire       [5:0]    _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2;
  wire       [5:0]    _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3;
  wire       [0:0]    _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3_1;
  wire       [5:0]    _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4;
  wire       [0:0]    _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4_1;
  wire       [5:0]    _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5;
  wire       [0:0]    _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5_1;
  wire       [5:0]    _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6;
  wire       [0:0]    _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6_1;
  wire       [11:0]   _zz__zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3;
  wire       [31:0]   _zz_ALU0_IntAluPlugin_logic_process_result;
  wire       [0:0]    _zz_ALU0_IntAluPlugin_logic_process_result_1;
  wire       [4:0]    _zz_ALU0_ShiftPlugin_logic_process_amplitude;
  wire       [31:0]   _zz_ALU0_ShiftPlugin_logic_process_reversed;
  wire                _zz_ALU0_ShiftPlugin_logic_process_reversed_1;
  wire       [0:0]    _zz_ALU0_ShiftPlugin_logic_process_reversed_2;
  wire       [20:0]   _zz_ALU0_ShiftPlugin_logic_process_reversed_3;
  wire                _zz_ALU0_ShiftPlugin_logic_process_reversed_4;
  wire       [0:0]    _zz_ALU0_ShiftPlugin_logic_process_reversed_5;
  wire       [9:0]    _zz_ALU0_ShiftPlugin_logic_process_reversed_6;
  wire       [32:0]   _zz_ALU0_ShiftPlugin_logic_process_shifted;
  wire       [32:0]   _zz_ALU0_ShiftPlugin_logic_process_shifted_1;
  wire       [31:0]   _zz_ALU0_ShiftPlugin_logic_process_patched;
  wire                _zz_ALU0_ShiftPlugin_logic_process_patched_1;
  wire       [0:0]    _zz_ALU0_ShiftPlugin_logic_process_patched_2;
  wire       [20:0]   _zz_ALU0_ShiftPlugin_logic_process_patched_3;
  wire                _zz_ALU0_ShiftPlugin_logic_process_patched_4;
  wire       [0:0]    _zz_ALU0_ShiftPlugin_logic_process_patched_5;
  wire       [9:0]    _zz_ALU0_ShiftPlugin_logic_process_patched_6;
  wire       [20:0]   _zz_ALU0_BranchPlugin_logic_process_target_b;
  wire       [11:0]   _zz_ALU0_BranchPlugin_logic_process_target_b_1;
  wire       [12:0]   _zz_ALU0_BranchPlugin_logic_process_target_b_2;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE;
  wire       [1:0]    _zz_ALU0_BranchPlugin_logic_process_slices;
  wire       [0:0]    _zz_ALU0_BranchPlugin_logic_process_slices_1;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE_1;
  wire       [11:0]   _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [11:0]   _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED_1;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED_1;
  wire       [46:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1;
  wire       [33:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_1;
  wire       [17:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_2;
  wire       [15:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_3;
  wire       [46:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2;
  wire       [33:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_1;
  wire       [15:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_2;
  wire       [17:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_3;
  wire       [29:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3;
  wire       [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3_1;
  wire       [15:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3_2;
  wire       [15:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3_3;
  wire       [62:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_3;
  wire       [62:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_4;
  wire       [62:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_5;
  wire       [62:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_6;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_3;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_4;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_5;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_6;
  wire       [34:0]   _zz_EU0_DivPlugin_logic_rsp_selected;
  wire       [34:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_1;
  wire       [34:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_2;
  wire       [34:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_3;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_4;
  wire       [11:0]   _zz__zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire       [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1;
  wire       [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3;
  wire       [31:0]   _zz_ALU1_IntAluPlugin_logic_process_result;
  wire       [0:0]    _zz_ALU1_IntAluPlugin_logic_process_result_1;
  wire       [4:0]    _zz_ALU1_ShiftPlugin_logic_process_amplitude;
  wire       [31:0]   _zz_ALU1_ShiftPlugin_logic_process_reversed;
  wire                _zz_ALU1_ShiftPlugin_logic_process_reversed_1;
  wire       [0:0]    _zz_ALU1_ShiftPlugin_logic_process_reversed_2;
  wire       [20:0]   _zz_ALU1_ShiftPlugin_logic_process_reversed_3;
  wire                _zz_ALU1_ShiftPlugin_logic_process_reversed_4;
  wire       [0:0]    _zz_ALU1_ShiftPlugin_logic_process_reversed_5;
  wire       [9:0]    _zz_ALU1_ShiftPlugin_logic_process_reversed_6;
  wire       [32:0]   _zz_ALU1_ShiftPlugin_logic_process_shifted;
  wire       [32:0]   _zz_ALU1_ShiftPlugin_logic_process_shifted_1;
  wire       [31:0]   _zz_ALU1_ShiftPlugin_logic_process_patched;
  wire                _zz_ALU1_ShiftPlugin_logic_process_patched_1;
  wire       [0:0]    _zz_ALU1_ShiftPlugin_logic_process_patched_2;
  wire       [20:0]   _zz_ALU1_ShiftPlugin_logic_process_patched_3;
  wire                _zz_ALU1_ShiftPlugin_logic_process_patched_4;
  wire       [0:0]    _zz_ALU1_ShiftPlugin_logic_process_patched_5;
  wire       [9:0]    _zz_ALU1_ShiftPlugin_logic_process_patched_6;
  wire       [20:0]   _zz_ALU1_BranchPlugin_logic_process_target_b;
  wire       [11:0]   _zz_ALU1_BranchPlugin_logic_process_target_b_1;
  wire       [12:0]   _zz_ALU1_BranchPlugin_logic_process_target_b_2;
  wire       [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TRUE;
  wire       [1:0]    _zz_ALU1_BranchPlugin_logic_process_slices;
  wire       [0:0]    _zz_ALU1_BranchPlugin_logic_process_slices_1;
  wire       [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE;
  wire       [3:0]    _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE_1;
  wire       [4:0]    _zz_BranchContextPlugin_logic_onCommit_commitedNext;
  reg        [1:0]    _zz_BranchContextPlugin_logic_onCommit_commitedNext_1;
  wire       [1:0]    _zz_BranchContextPlugin_logic_onCommit_commitedNext_2;
  wire       [24:0]   _zz_HistoryPlugin_logic_onCommit_valueNext_1;
  wire       [24:0]   _zz_HistoryPlugin_logic_onCommit_valueNext_2;
  wire       [24:0]   _zz_HistoryPlugin_logic_update_pushes_0_stateNext_1;
  wire       [24:0]   _zz_HistoryPlugin_logic_update_pushes_2_stateNext_1;
  wire       [24:0]   _zz_HistoryPlugin_logic_update_pushes_2_stateNext_2;
  reg        [23:0]   _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_2;
  wire       [0:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_3;
  reg        [0:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_2;
  wire       [0:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_3;
  wire       [0:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken;
  wire       [0:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken_1;
  reg        [3:0]    _zz_DecoderPredictionPlugin_logic_ras_healPush_2;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_ras_healPush_3;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_tracker_freeNext;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_tracker_freeNext_1;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_tracker_freeNext_2;
  reg        [1:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount;
  wire       [1:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount_1;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_1;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_2;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_3;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_4;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_5;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_6;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_7;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_8;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_9;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_10;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_11;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_12;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_13;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_14;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_15;
  wire       [14:0]   _zz_Lsu2Plugin_logic_lq_onCommit_priority_1;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_onCommit_free_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_onCommit_free_1_1;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_16;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_17;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_18;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_19;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_20;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_21;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_22;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_23;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_24;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_25;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_26;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_27;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_28;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_29;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_30;
  wire       [3:0]    _zz_when_Lsu2Plugin_l454_31;
  wire       [14:0]   _zz_Lsu2Plugin_logic_lq_onCommit_priority_2;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_onCommit_free_2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_onCommit_free_2_1;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_ptr_free;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext_1;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext_2;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext_3;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeNext_4;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1_1;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_2_1;
  reg        [1:0]    _zz_Lsu2Plugin_logic_allocation_loads_requestsCount;
  wire       [1:0]    _zz_Lsu2Plugin_logic_allocation_loads_requestsCount_1;
  reg        [1:0]    _zz_Lsu2Plugin_logic_allocation_stores_requestsCount;
  wire       [1:0]    _zz_Lsu2Plugin_logic_allocation_stores_requestsCount_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_spFpAddress_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_spFpAddress_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_addressPre_port;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_addressPre_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_physRd_port;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_physRd_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_robId_port;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_robId_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_pc_port;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_pc_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_writeRd_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_writeRd_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_lr_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_lr_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_size_port;
  wire       [1:0]    _zz_Lsu2Plugin_logic_lq_mem_size_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_unsigned_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_unsigned_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port;
  wire       [2:0]    _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port;
  wire       [5:0]    _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_addressPre_port;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_addressPre_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_robId_port;
  wire       [5:0]    _zz_Lsu2Plugin_logic_sq_mem_robId_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_amo_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_amo_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_sc_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_sc_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_size_port;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sq_mem_size_port_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_data_port;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_1;
  wire       [15:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh;
  wire       [15:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh;
  wire       [6:0]    _zz_Lsu2Plugin_logic_lqSqArbitration_s1_cmp;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu_1;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_1;
  wire       [4:0]    _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT;
  wire       [4:0]    _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_3;
  wire       [7:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_4;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_5;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_6;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_3;
  wire       [7:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_4;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_5;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_6;
  wire                _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input_2;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input_3;
  wire                _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits_2;
  wire       [5:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits_3;
  wire       [15:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh_1;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh_2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_lq_mem_addressPost_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_lq_mem_io_port;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sq_mem_addressPost_port;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_mem_io_port;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_3;
  wire       [7:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_4;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_5;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_6;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_3;
  wire       [7:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_4;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_5;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_6;
  wire       [15:0]   _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh;
  reg        [7:0]    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_1;
  reg        [7:0]    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_2;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_3;
  reg                 _zz__zz_when_Lsu2Plugin_l1348;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_1;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_2;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_1;
  wire       [6:0]    _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_2;
  wire       [1:0]    _zz_when_SInt_l132;
  wire       [0:0]    _zz_when_SInt_l138;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sq_ptr_writeBack;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sq_ptr_writeBack_1;
  wire       [2:0]    _zz_Lsu2Plugin_setup_specialTrap_payload_cause;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_3;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_4;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_5;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_6;
  wire       [1:0]    _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_7;
  wire       [31:0]   _zz_ALU0_BranchPlugin_setup_intFormatPort_payload;
  wire       [4:0]    _zz_ALU0_BranchPlugin_setup_reschedule_payload_reason;
  wire       [31:0]   _zz_ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice;
  wire       [1:0]    _zz_ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice_1;
  wire       [31:0]   _zz_ALU1_BranchPlugin_setup_intFormatPort_payload;
  wire       [4:0]    _zz_ALU1_BranchPlugin_setup_reschedule_payload_reason;
  wire       [31:0]   _zz_ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice;
  wire       [1:0]    _zz_ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice_1;
  wire       [41:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port_1;
  wire       [41:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port_1;
  wire       [41:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port_1;
  wire       [41:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port_1;
  wire       [1:0]    _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
  wire       [0:0]    _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1;
  wire       [21:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port_1;
  wire       [21:0]   _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port_1;
  wire       [41:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port_1;
  wire       [41:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port_1;
  wire       [41:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port_1;
  wire       [41:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port_1;
  wire       [1:0]    _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
  wire       [0:0]    _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1;
  wire       [21:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port_1;
  wire       [21:0]   _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port_1;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_6;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_1;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_2;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_3;
  wire       [11:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_4;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_5;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_6;
  wire       [11:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_7;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_8;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_9;
  wire       [11:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_10;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_11;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_12;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_13;
  wire       [0:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault;
  wire       [4:0]    _zz_PerformanceCounterPlugin_setup_readPort_address;
  wire       [4:0]    _zz_PerformanceCounterPlugin_setup_writePort_address;
  wire       [58:0]   _zz_PerformanceCounterPlugin_logic_fsm_calc;
  wire       [58:0]   _zz_PerformanceCounterPlugin_logic_fsm_calc_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_fsm_calc_2;
  wire       [4:0]    _zz_PerformanceCounterPlugin_logic_fsm_calc_3;
  wire       [6:0]    _zz_PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_6;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineException;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_1;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_2;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_3;
  wire       [11:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_4;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_5;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_6;
  wire       [11:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_7;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_8;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_9;
  wire       [11:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_10;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_11;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_12;
  wire       [31:0]   _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_13;
  wire       [0:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault;
  wire       [1:0]    _zz_MmuPlugin_logic_refill_portsRequests_ohFirst_masked;
  wire       [3:0]    _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask_1;
  wire       [3:0]    _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask_1;
  wire       [1:0]    _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask;
  wire       [1:0]    _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask;
  wire       [3:0]    _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  reg        [4:0]    _zz_CsrRamPlugin_logic_writeLogic_port_payload_address;
  reg        [31:0]   _zz_CsrRamPlugin_logic_writeLogic_port_payload_data;
  wire       [2:0]    _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  reg        [4:0]    _zz_CsrRamPlugin_logic_readLogic_port_address;
  wire       [11:0]   _zz_COMB_CSR_;
  wire       [11:0]   _zz_COMB_CSR__1;
  wire                _zz_COMB_CSR__2;
  wire       [0:0]    _zz_COMB_CSR__3;
  wire       [79:0]   _zz_COMB_CSR__4;
  wire       [11:0]   _zz_COMB_CSR__5;
  wire       [11:0]   _zz_COMB_CSR__6;
  wire                _zz_COMB_CSR__7;
  wire       [0:0]    _zz_COMB_CSR__8;
  wire       [72:0]   _zz_COMB_CSR__9;
  wire       [11:0]   _zz_COMB_CSR__10;
  wire       [11:0]   _zz_COMB_CSR__11;
  wire                _zz_COMB_CSR__12;
  wire       [0:0]    _zz_COMB_CSR__13;
  wire       [65:0]   _zz_COMB_CSR__14;
  wire       [11:0]   _zz_COMB_CSR__15;
  wire       [11:0]   _zz_COMB_CSR__16;
  wire                _zz_COMB_CSR__17;
  wire       [0:0]    _zz_COMB_CSR__18;
  wire       [58:0]   _zz_COMB_CSR__19;
  wire       [11:0]   _zz_COMB_CSR__20;
  wire       [11:0]   _zz_COMB_CSR__21;
  wire                _zz_COMB_CSR__22;
  wire       [0:0]    _zz_COMB_CSR__23;
  wire       [51:0]   _zz_COMB_CSR__24;
  wire       [11:0]   _zz_COMB_CSR__25;
  wire       [11:0]   _zz_COMB_CSR__26;
  wire                _zz_COMB_CSR__27;
  wire       [0:0]    _zz_COMB_CSR__28;
  wire       [44:0]   _zz_COMB_CSR__29;
  wire       [11:0]   _zz_COMB_CSR__30;
  wire       [11:0]   _zz_COMB_CSR__31;
  wire                _zz_COMB_CSR__32;
  wire       [0:0]    _zz_COMB_CSR__33;
  wire       [37:0]   _zz_COMB_CSR__34;
  wire       [11:0]   _zz_COMB_CSR__35;
  wire       [11:0]   _zz_COMB_CSR__36;
  wire                _zz_COMB_CSR__37;
  wire       [0:0]    _zz_COMB_CSR__38;
  wire       [30:0]   _zz_COMB_CSR__39;
  wire       [11:0]   _zz_COMB_CSR__40;
  wire       [11:0]   _zz_COMB_CSR__41;
  wire                _zz_COMB_CSR__42;
  wire       [0:0]    _zz_COMB_CSR__43;
  wire       [23:0]   _zz_COMB_CSR__44;
  wire       [11:0]   _zz_COMB_CSR__45;
  wire       [11:0]   _zz_COMB_CSR__46;
  wire                _zz_COMB_CSR__47;
  wire       [0:0]    _zz_COMB_CSR__48;
  wire       [16:0]   _zz_COMB_CSR__49;
  wire       [11:0]   _zz_COMB_CSR__50;
  wire       [11:0]   _zz_COMB_CSR__51;
  wire                _zz_COMB_CSR__52;
  wire       [0:0]    _zz_COMB_CSR__53;
  wire       [9:0]    _zz_COMB_CSR__54;
  wire       [11:0]   _zz_COMB_CSR__55;
  wire       [11:0]   _zz_COMB_CSR__56;
  wire                _zz_COMB_CSR__57;
  wire       [0:0]    _zz_COMB_CSR__58;
  wire       [2:0]    _zz_COMB_CSR__59;
  wire       [11:0]   _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter;
  wire       [11:0]   _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_1;
  wire                _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_2;
  wire       [0:0]    _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_3;
  wire       [16:0]   _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_4;
  wire       [11:0]   _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_5;
  wire       [11:0]   _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_6;
  wire                _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_7;
  wire       [0:0]    _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_8;
  wire       [9:0]    _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_9;
  wire       [11:0]   _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_10;
  wire       [11:0]   _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_11;
  wire                _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_12;
  wire       [0:0]    _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_13;
  wire       [2:0]    _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_14;
  wire       [0:0]    _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented;
  wire       [21:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_1;
  wire       [0:0]    _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_2;
  wire       [10:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_3;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_setup_onDecodeAddress;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_setup_onReadAddress;
  reg        [31:0]   _zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17;
  wire       [0:0]    _zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17_1;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [4:0]    _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_setup_onWriteAddress;
  wire       [31:0]   _zz_csrAccess_payload_address;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_2;
  wire                _zz_FrontendPlugin_decoded_LEGAL_0_3;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_4;
  wire       [18:0]   _zz_FrontendPlugin_decoded_LEGAL_0_5;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_6;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_7;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_8;
  wire                _zz_FrontendPlugin_decoded_LEGAL_0_9;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_10;
  wire       [12:0]   _zz_FrontendPlugin_decoded_LEGAL_0_11;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_12;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_13;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_14;
  wire                _zz_FrontendPlugin_decoded_LEGAL_0_15;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_16;
  wire       [6:0]    _zz_FrontendPlugin_decoded_LEGAL_0_17;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_18;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_19;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_0_20;
  wire                _zz_FrontendPlugin_decoded_LEGAL_0_21;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_22;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_0_23;
  wire       [0:0]    _zz_FrontendPlugin_decoded_READ_RS_0_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_READ_RS_1_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_WRITE_RD_0_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_WRITE_RD_0_2;
  wire       [31:0]   _zz_FrontendPlugin_decoded_WRITE_RD_0_3;
  wire       [31:0]   _zz_FrontendPlugin_decoded_WRITE_RD_0_4;
  wire                _zz_FrontendPlugin_decoded_WRITE_RD_0_5;
  wire       [0:0]    _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_0_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_EU0_SEL_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LQ_ALLOC_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_SQ_ALLOC_0_2;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_2;
  wire                _zz_FrontendPlugin_decoded_LEGAL_1_3;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_1_4;
  wire       [18:0]   _zz_FrontendPlugin_decoded_LEGAL_1_5;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_6;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_7;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_8;
  wire                _zz_FrontendPlugin_decoded_LEGAL_1_9;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_1_10;
  wire       [12:0]   _zz_FrontendPlugin_decoded_LEGAL_1_11;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_12;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_13;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_14;
  wire                _zz_FrontendPlugin_decoded_LEGAL_1_15;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_1_16;
  wire       [6:0]    _zz_FrontendPlugin_decoded_LEGAL_1_17;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_18;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_19;
  wire       [31:0]   _zz_FrontendPlugin_decoded_LEGAL_1_20;
  wire                _zz_FrontendPlugin_decoded_LEGAL_1_21;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_1_22;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LEGAL_1_23;
  wire       [0:0]    _zz_FrontendPlugin_decoded_READ_RS_0_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_READ_RS_1_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_WRITE_RD_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_WRITE_RD_1_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_WRITE_RD_1_2;
  wire       [31:0]   _zz_FrontendPlugin_decoded_WRITE_RD_1_3;
  wire                _zz_FrontendPlugin_decoded_WRITE_RD_1_4;
  wire       [0:0]    _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_1_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_EU0_SEL_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_LQ_ALLOC_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_SQ_ALLOC_1_2;
  wire       [1:0]    _zz__zz_DecoderPlugin_setup_exceptionPort_payload_tval_1;
  wire       [1:0]    _zz__zz_DecoderPlugin_setup_exceptionPort_payload_tval_1_1;
  wire       [0:0]    _zz_DecoderPlugin_logic_exception_fetchFault;
  wire       [0:0]    _zz_DecoderPlugin_logic_exception_fetchFaultPage;
  wire       [0:0]    _zz_DecoderPlugin_logic_exception_debugEnter;
  wire       [31:0]   _zz_DecoderPlugin_setup_exceptionPort_payload_tval_2;
  wire       [31:0]   _zz_DecoderPlugin_setup_exceptionPort_payload_tval_3;
  wire       [1:0]    _zz_DecoderPlugin_setup_exceptionPort_payload_tval_4;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_2;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_3;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_2;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_3;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_2;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_3;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_2;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_3;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_1_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_1_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_1;
  wire       [0:0]    _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_1_1;
  wire       [11:0]   _zz_FrontendPlugin_decoded_OP_ID;
  wire       [1:0]    _zz_FrontendPlugin_decoded_OP_ID_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_IS_JAL_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_IS_JALR_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_Prediction_IS_BRANCH_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_IS_ANY_0_1;
  wire       [12:0]   _zz__zz_FrontendPlugin_decoded_OFFSET_0;
  wire       [20:0]   _zz__zz_FrontendPlugin_decoded_OFFSET_0_1;
  wire       [1:0]    _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_PC_INC_0;
  wire       [31:0]   _zz_FrontendPlugin_decoded_PC_INC_0_1;
  wire       [3:0]    _zz_FrontendPlugin_decoded_PC_INC_0_2;
  wire       [31:0]   _zz_FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0;
  wire       [0:0]    _zz_FrontendPlugin_decoded_IS_JAL_1_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_IS_JALR_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_Prediction_IS_BRANCH_1;
  wire       [0:0]    _zz_FrontendPlugin_decoded_IS_ANY_1_1;
  wire       [12:0]   _zz__zz_FrontendPlugin_decoded_OFFSET_1;
  wire       [20:0]   _zz__zz_FrontendPlugin_decoded_OFFSET_1_1;
  wire       [1:0]    _zz_DecoderPredictionPlugin_logic_decodePatch_slots_1_pcAdd_slices;
  wire       [0:0]    _zz_DecoderPredictionPlugin_logic_decodePatch_slots_1_pcAdd_slices_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_PC_INC_1;
  wire       [31:0]   _zz_FrontendPlugin_decoded_PC_INC_1_1;
  wire       [3:0]    _zz_FrontendPlugin_decoded_PC_INC_1_2;
  wire       [31:0]   _zz_FrontendPlugin_decoded_PC_TARGET_PRE_RAS_1;
  wire       [31:0]   _zz_DecoderPredictionPlugin_setup_decodeJump_payload_pc;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2;
  wire       [5:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_1;
  wire       [5:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2;
  wire       [5:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_1;
  wire       [5:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_1;
  wire       [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_2;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_1;
  wire       [3:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_2;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
  wire       [0:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1;
  wire       [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1;
  wire       [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2;
  wire       [5:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_1;
  wire       [5:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_2;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2;
  wire       [5:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_1;
  wire       [5:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_2;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2;
  wire       [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PC_1;
  wire       [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PC_2;
  wire       [3:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_1;
  wire       [3:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_2;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_2;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_2;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
  wire       [0:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_3;
  reg        [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_3;
  reg        [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_3;
  reg        [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_3;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_3;
  reg        [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_3;
  reg        [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_3;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_2;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire       [0:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1;
  wire                _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0;
  wire       [0:0]    _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_1;
  wire       [22:0]   _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_2;
  wire                _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_3;
  wire       [0:0]    _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_4;
  wire       [14:0]   _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_5;
  wire                _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_6;
  wire       [0:0]    _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_7;
  wire       [6:0]    _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_8;
  wire       [5:0]    _zz_DispatchPlugin_logic_ptr_next;
  wire       [4:0]    _zz_DispatchPlugin_logic_push_commitNotWaitingOnUs;
  wire       [31:0]   _zz_DispatchPlugin_logic_push_slots_0_events_0;
  wire       [4:0]    _zz_DispatchPlugin_logic_push_slots_0_events_0_1;
  wire       [5:0]    _zz_DispatchPlugin_logic_push_slots_0_events_0_2;
  wire       [31:0]   _zz_DispatchPlugin_logic_push_slots_0_events_1;
  wire       [4:0]    _zz_DispatchPlugin_logic_push_slots_0_events_1_1;
  wire       [5:0]    _zz_DispatchPlugin_logic_push_slots_0_events_1_2;
  wire       [31:0]   _zz_DispatchPlugin_logic_push_slots_1_events_0;
  wire       [4:0]    _zz_DispatchPlugin_logic_push_slots_1_events_0_1;
  wire       [5:0]    _zz_DispatchPlugin_logic_push_slots_1_events_0_2;
  wire       [31:0]   _zz_DispatchPlugin_logic_push_slots_1_events_1;
  wire       [4:0]    _zz_DispatchPlugin_logic_push_slots_1_events_1_1;
  wire       [5:0]    _zz_DispatchPlugin_logic_push_slots_1_events_1_2;
  wire                _zz_DispatchPlugin_logic_pop_0_portEventFull;
  wire       [0:0]    _zz_DispatchPlugin_logic_pop_0_portEventFull_1;
  wire       [21:0]   _zz_DispatchPlugin_logic_pop_0_portEventFull_2;
  wire                _zz_DispatchPlugin_logic_pop_0_portEventFull_3;
  wire       [0:0]    _zz_DispatchPlugin_logic_pop_0_portEventFull_4;
  wire       [10:0]   _zz_DispatchPlugin_logic_pop_0_portEventFull_5;
  wire                _zz_DispatchPlugin_logic_pop_0_portEventFull_6;
  wire                _zz_DispatchPlugin_logic_pop_0_portEventFull_7;
  wire       [5:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID;
  wire                _zz_DispatchPlugin_logic_pop_1_portEventFull;
  wire       [0:0]    _zz_DispatchPlugin_logic_pop_1_portEventFull_1;
  wire       [21:0]   _zz_DispatchPlugin_logic_pop_1_portEventFull_2;
  wire                _zz_DispatchPlugin_logic_pop_1_portEventFull_3;
  wire       [0:0]    _zz_DispatchPlugin_logic_pop_1_portEventFull_4;
  wire       [12:0]   _zz_DispatchPlugin_logic_pop_1_portEventFull_5;
  wire                _zz_DispatchPlugin_logic_pop_1_portEventFull_6;
  wire       [0:0]    _zz_DispatchPlugin_logic_pop_1_portEventFull_7;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_1_portEventFull_8;
  wire       [5:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID;
  wire                _zz_DispatchPlugin_logic_pop_2_portEventFull;
  wire       [0:0]    _zz_DispatchPlugin_logic_pop_2_portEventFull_1;
  wire       [22:0]   _zz_DispatchPlugin_logic_pop_2_portEventFull_2;
  wire                _zz_DispatchPlugin_logic_pop_2_portEventFull_3;
  wire       [0:0]    _zz_DispatchPlugin_logic_pop_2_portEventFull_4;
  wire       [11:0]   _zz_DispatchPlugin_logic_pop_2_portEventFull_5;
  wire                _zz_DispatchPlugin_logic_pop_2_portEventFull_6;
  wire       [0:0]    _zz_DispatchPlugin_logic_pop_2_portEventFull_7;
  wire       [0:0]    _zz_DispatchPlugin_logic_pop_2_portEventFull_8;
  wire       [5:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_1_ROB_ID;
  wire       [5:0]    _zz_DispatchPlugin_logic_wake_dynamic_offseted_0_payload;
  wire       [5:0]    _zz_DispatchPlugin_logic_wake_dynamic_offseted_1_payload;
  wire       [5:0]    _zz_DispatchPlugin_logic_wake_dynamic_offseted_2_payload;
  wire       [5:0]    _zz_DispatchPlugin_logic_wake_dynamic_offseted_3_payload;
  wire       [31:0]   _zz_DispatchPlugin_logic_wake_dynamic_masks_0;
  wire       [31:0]   _zz_DispatchPlugin_logic_wake_dynamic_masks_1;
  wire       [31:0]   _zz_DispatchPlugin_logic_wake_dynamic_masks_2;
  wire       [31:0]   _zz_DispatchPlugin_logic_wake_dynamic_masks_3;
  reg        [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_3;
  reg        [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_3;
  reg        [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_3;
  reg        [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_3;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_3;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_3;
  wire       [4:0]    _zz_RobPlugin_logic_completionMem_init_0_robId;
  wire       [4:0]    _zz_RobPlugin_logic_completionMem_init_1_robId;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_0_port;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_1_port;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_2_port;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_3_port;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_4_port;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_5_port;
  wire       [0:0]    _zz_RobPlugin_logic_completionMem_hits_6_port;
  wire       [4:0]    _zz__zz_CommitPlugin_setup_robLineMask_mask;
  wire       [4:0]    _zz__zz_CommitPlugin_setup_robLineMask_mask_1;
  wire       [4:0]    _zz__zz_when_RobPlugin_l118;
  wire       [4:0]    _zz__zz_when_RobPlugin_l118_1;
  wire       [4:0]    _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port;
  wire       [1:0]    _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port_1;
  wire                _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port_2;
  wire       [1:0]    _zz__zz_CommitPlugin_logic_commit_active_2;
  wire       [1:0]    _zz__zz_integer_RfAllocationPlugin_logic_push_mask_0_2;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_PC_banks_0_port_1;
  wire       [31:0]   _zz_RobPlugin_logic_storage_PC_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_PC_banks_1_port_1;
  wire       [63:0]   _zz__zz_commit_pc_0_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port_1;
  wire       [1:0]    _zz__zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1;
  wire       [1:0]    _zz__zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1;
  wire       [4:0]    _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port;
  wire       [11:0]   _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port_1;
  wire                _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port_2;
  wire       [11:0]   _zz__zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2;
  wire       [11:0]   _zz__zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2;
  wire       [4:0]    _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port;
  wire       [9:0]    _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port_1;
  wire                _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port_2;
  wire       [9:0]    _zz__zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2;
  wire       [4:0]    _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port;
  wire       [11:0]   _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port_1;
  wire                _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port_2;
  wire       [11:0]   _zz__zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2;
  wire       [4:0]    _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port;
  wire       [1:0]    _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port_1;
  wire                _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port_2;
  wire       [1:0]    _zz__zz_BranchContextPlugin_logic_onCommit_isBranch_0_2;
  wire       [0:0]    _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port_1;
  wire       [1:0]    _zz__zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1;
  wire                _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_1_port;
  wire       [3:0]    _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port_1;
  wire       [3:0]    _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1_port_1;
  wire       [4:0]    _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port;
  wire       [1:0]    _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port_1;
  wire                _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port_2;
  wire       [1:0]    _zz__zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2;
  wire       [4:0]    _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port;
  wire       [1:0]    _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port_1;
  wire                _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port_2;
  wire       [1:0]    _zz__zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2;
  wire                _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1_port;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port_1;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_1_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port_1;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port_1;
  wire       [5:0]    _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_1_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port_1;
  wire       [3:0]    _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port_1;
  wire       [3:0]    _zz_RobPlugin_logic_storage_BRANCH_ID_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_BRANCH_ID_banks_1_port_1;
  wire       [4:0]    _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port_1;
  wire       [4:0]    _zz_RobPlugin_logic_storage_LSU_ID_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_LSU_ID_banks_1_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port;
  wire                _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port_1;
  wire       [0:0]    _zz_RobPlugin_logic_storage_ROB_MSB_banks_1_port;
  wire                _zz_RobPlugin_logic_storage_ROB_MSB_banks_1_port_1;
  wire       [6:0]    _zz_PcPlugin_logic_init_counter;
  wire       [0:0]    _zz_PcPlugin_logic_init_counter_1;
  wire       [31:0]   _zz_PcPlugin_logic_fetchPc_pc;
  wire       [3:0]    _zz_PcPlugin_logic_fetchPc_pc_1;
  reg        [5:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_11;
  wire       [63:0]   _zz_PerformanceCounterPlugin_setup_writePort_data;
  wire       [31:0]   _zz_PerformanceCounterPlugin_setup_writePort_data_1;
  wire       [4:0]    _zz_PerformanceCounterPlugin_setup_writePort_address_1;
  wire       [31:0]   _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded;
  wire       [31:0]   _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2_1;
  wire       [31:0]   _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3_2;
  wire       [31:0]   _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4_2;
  wire       [31:0]   _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5_2;
  wire       [31:0]   _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6_2;
  wire       [31:0]   _zz_PrivilegedPlugin_setup_ramWrite_data;
  wire       [31:0]   _zz_PrivilegedPlugin_setup_ramWrite_data_1;
  wire       [31:0]   _zz_PrivilegedPlugin_logic_readed;
  wire       [31:0]   _zz_PrivilegedPlugin_logic_readed_1;
  wire       [3:0]    _zz_PrivilegedPlugin_logic_readed_2;
  wire       [3:0]    _zz_PrivilegedPlugin_logic_readed_3;
  wire       [1:0]    _zz_PrivilegedPlugin_logic_readed_4;
  wire       [1:0]    _zz_PrivilegedPlugin_logic_readed_5;
  wire       [0:0]    _zz_PrivilegedPlugin_logic_readed_6;
  wire                FetchPlugin_stages_2_isFlushingRoot;
  wire                FetchPlugin_stages_1_isFlushingRoot;
  wire                FetchPlugin_stages_0_isFlushed;
  wire                FetchPlugin_stages_1_isFlushingNext;
  wire                FetchPlugin_stages_1_isThrown;
  wire                FetchPlugin_stages_2_isFlushed;
  reg        [31:0]   FetchPlugin_stages_2_Fetch_FETCH_PC_INC;
  reg        [1:0]    FetchPlugin_stages_2_GSHARE_COUNTER_0;
  reg        [1:0]    FetchPlugin_stages_2_GSHARE_COUNTER_1;
  reg                 FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE;
  reg        [0:0]    FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_SLICE;
  reg                 FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID;
  reg        [31:0]   FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT;
  reg        [1:0]    FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT;
  reg                 FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID;
  reg        [0:0]    FetchPlugin_stages_2_Prediction_WORD_BRANCH_SLICE;
  reg        [23:0]   FetchPlugin_stages_1_BRANCH_HISTORY;
  reg        [11:0]   FetchPlugin_stages_2_FETCH_ID;
  reg        [31:0]   FetchPlugin_stages_1_Fetch_FETCH_PC_INC;
  wire                FrontendPlugin_dispatch_isFlushingRoot;
  wire                FrontendPlugin_decoded_isFlushingRoot;
  wire                FrontendPlugin_decompressed_isFlushed;
  wire                FrontendPlugin_allocated_isFlushed;
  wire                FrontendPlugin_dispatch_isFlushed;
  wire                FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_1_1;
  wire                FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_0_1;
  wire                FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_1_0;
  wire                FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_0_0;
  wire                FrontendPlugin_allocated_EU0_SEL_1;
  reg                 FrontendPlugin_serialized_EU0_SEL_1;
  wire                FrontendPlugin_allocated_ALU0_ALU1_SEL_1;
  reg                 FrontendPlugin_serialized_ALU0_ALU1_SEL_1;
  wire                FrontendPlugin_allocated_EU0_SEL_0;
  reg                 FrontendPlugin_serialized_EU0_SEL_0;
  wire                FrontendPlugin_allocated_ALU0_ALU1_SEL_0;
  reg                 FrontendPlugin_serialized_ALU0_ALU1_SEL_0;
  wire                FrontendPlugin_allocated_DispatchPlugin_FENCE_YOUNGER_1;
  wire                FrontendPlugin_allocated_DispatchPlugin_FENCE_YOUNGER_0;
  wire                FrontendPlugin_allocated_DispatchPlugin_FENCE_OLDER_1;
  wire                FrontendPlugin_allocated_DispatchPlugin_FENCE_OLDER_0;
  wire       [1:0]    FrontendPlugin_allocated_GSHARE_COUNTER_1_0;
  wire       [1:0]    FrontendPlugin_allocated_GSHARE_COUNTER_1_1;
  reg        [1:0]    FrontendPlugin_serialized_GSHARE_COUNTER_1_0;
  reg        [1:0]    FrontendPlugin_serialized_GSHARE_COUNTER_1_1;
  wire       [1:0]    FrontendPlugin_decoded_GSHARE_COUNTER_1_0;
  wire       [1:0]    FrontendPlugin_decoded_GSHARE_COUNTER_1_1;
  wire       [1:0]    FrontendPlugin_allocated_GSHARE_COUNTER_0_0;
  wire       [1:0]    FrontendPlugin_allocated_GSHARE_COUNTER_0_1;
  reg        [1:0]    FrontendPlugin_serialized_GSHARE_COUNTER_0_0;
  reg        [1:0]    FrontendPlugin_serialized_GSHARE_COUNTER_0_1;
  wire       [1:0]    FrontendPlugin_decoded_GSHARE_COUNTER_0_0;
  wire       [1:0]    FrontendPlugin_decoded_GSHARE_COUNTER_0_1;
  wire                FrontendPlugin_allocated_Prediction_IS_BRANCH_1;
  wire                FrontendPlugin_allocated_Prediction_IS_BRANCH_0;
  wire                FrontendPlugin_allocated_SQ_ALLOC_1;
  reg                 FrontendPlugin_serialized_SQ_ALLOC_1;
  wire                FrontendPlugin_allocated_SQ_ALLOC_0;
  reg                 FrontendPlugin_serialized_SQ_ALLOC_0;
  wire                FrontendPlugin_allocated_LQ_ALLOC_1;
  reg                 FrontendPlugin_serialized_LQ_ALLOC_1;
  wire                FrontendPlugin_allocated_LQ_ALLOC_0;
  reg                 FrontendPlugin_serialized_LQ_ALLOC_0;
  reg        [11:0]   FrontendPlugin_serialized_OP_ID;
  reg        [23:0]   FrontendPlugin_serialized_BRANCH_HISTORY_1;
  wire       [23:0]   FrontendPlugin_decoded_BRANCH_HISTORY_1;
  wire       [23:0]   FrontendPlugin_decompressed_BRANCH_HISTORY_1;
  reg        [23:0]   FrontendPlugin_serialized_BRANCH_HISTORY_0;
  wire       [23:0]   FrontendPlugin_decoded_BRANCH_HISTORY_0;
  wire       [23:0]   FrontendPlugin_decompressed_BRANCH_HISTORY_0;
  reg                 FrontendPlugin_serialized_READ_RS_1_1;
  reg        [4:0]    FrontendPlugin_serialized_ARCH_RS_1_1;
  reg                 FrontendPlugin_serialized_READ_RS_0_1;
  reg        [4:0]    FrontendPlugin_serialized_ARCH_RS_0_1;
  reg                 FrontendPlugin_serialized_READ_RS_1_0;
  reg        [4:0]    FrontendPlugin_serialized_ARCH_RS_1_0;
  reg                 FrontendPlugin_serialized_READ_RS_0_0;
  reg        [4:0]    FrontendPlugin_serialized_ARCH_RS_0_0;
  reg        [4:0]    FrontendPlugin_serialized_ARCH_RD_1;
  reg        [4:0]    FrontendPlugin_serialized_ARCH_RD_0;
  reg        [31:0]   FrontendPlugin_serialized_PC_1;
  reg        [31:0]   FrontendPlugin_serialized_PC_0;
  reg                 FrontendPlugin_serialized_WRITE_RD_1;
  reg                 FrontendPlugin_serialized_WRITE_RD_0;
  reg        [11:0]   FrontendPlugin_serialized_FETCH_ID_1;
  reg        [11:0]   FrontendPlugin_serialized_FETCH_ID_0;
  wire                FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_VALID_1;
  wire                FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_VALID_1;
  wire                FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_VALID_0;
  wire                FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_VALID_0;
  wire       [31:0]   FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_PC_NEXT_1;
  wire       [31:0]   FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  wire       [31:0]   FrontendPlugin_decompressed_PC_1;
  wire       [31:0]   FrontendPlugin_decompressed_PC_0;
  wire                FrontendPlugin_decompressed_Frontend_FETCH_FAULT_PAGE_1;
  wire                FrontendPlugin_decompressed_Frontend_FETCH_FAULT_PAGE_0;
  wire                FrontendPlugin_decompressed_Frontend_FETCH_FAULT_1;
  wire                FrontendPlugin_decompressed_Frontend_MASK_ALIGNED_1;
  wire                FrontendPlugin_decompressed_Frontend_FETCH_FAULT_0;
  wire                FrontendPlugin_decompressed_Frontend_MASK_ALIGNED_0;
  wire       [11:0]   FrontendPlugin_decompressed_FETCH_ID_1;
  wire       [11:0]   FrontendPlugin_decompressed_FETCH_ID_0;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_1_1;
  reg        [4:0]    FrontendPlugin_dispatch_ARCH_RS_1_1;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1;
  reg                 FrontendPlugin_dispatch_READ_RS_1_1;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_0_1;
  reg        [4:0]    FrontendPlugin_dispatch_ARCH_RD_0;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1;
  reg                 FrontendPlugin_dispatch_READ_RS_0_1;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_1_0;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0;
  reg                 FrontendPlugin_dispatch_READ_RS_1_0;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_0_0;
  reg                 FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0;
  reg                 FrontendPlugin_dispatch_READ_RS_0_0;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 _zz_3;
  reg                 _zz_4;
  reg                 _zz_5;
  reg                 _zz_6;
  reg                 _zz_7;
  reg                 _zz_8;
  wire                DispatchPlugin_logic_pop_2_stagesList_0_isFlushed;
  wire                DispatchPlugin_logic_pop_2_stagesList_1_isFlushed;
  reg                 DispatchPlugin_logic_pop_2_stagesList_1_ready;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_0;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_1;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_2;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_3;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_4;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_5;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_6;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_7;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_8;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_9;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_10;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_PHYS_RS_1;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_0;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_1;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_2;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_3;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_4;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_5;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_6;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_7;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_8;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_9;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_10;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_0;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_1;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_2;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_3;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_4;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_5;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_6;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_7;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_8;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_9;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_10;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_PHYS_RS_0;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_0;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_1;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_2;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_3;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_4;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_5;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_6;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_7;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_8;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_9;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_10;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_0;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_1;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_2;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_3;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_4;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_5;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_6;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_7;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_8;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_9;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_10;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_PHYS_RD;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_0;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_1;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_2;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_3;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_4;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_5;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_6;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_7;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_8;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_9;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_10;
  wire                DispatchPlugin_logic_pop_2_stagesList_0_LATENCY_0;
  reg        [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_OFFSET;
  reg        [4:0]    DispatchPlugin_logic_pop_2_stagesList_1_UINT;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_1_ROB_ID;
  wire       [4:0]    DispatchPlugin_logic_pop_2_stagesList_0_UINT;
  wire                DispatchPlugin_logic_pop_2_stagesList_0_ready;
  wire       [5:0]    DispatchPlugin_logic_pop_2_stagesList_0_OFFSET;
  wire       [31:0]   DispatchPlugin_logic_pop_2_stagesList_0_OH;
  wire                DispatchPlugin_logic_pop_1_stagesList_0_isFlushed;
  wire                DispatchPlugin_logic_pop_1_stagesList_1_isFlushed;
  reg                 DispatchPlugin_logic_pop_1_stagesList_1_LATENCY_0;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_0;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_1;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_2;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_3;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_4;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_5;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RD;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_0;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_1;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_2;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_3;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_4;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_5;
  wire                DispatchPlugin_logic_pop_1_stagesList_0_LATENCY_0;
  reg        [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_OFFSET;
  reg        [4:0]    DispatchPlugin_logic_pop_1_stagesList_1_UINT;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID;
  wire       [4:0]    DispatchPlugin_logic_pop_1_stagesList_0_UINT;
  wire                DispatchPlugin_logic_pop_1_stagesList_0_ready;
  wire       [5:0]    DispatchPlugin_logic_pop_1_stagesList_0_OFFSET;
  wire       [31:0]   DispatchPlugin_logic_pop_1_stagesList_0_OH;
  wire                DispatchPlugin_logic_pop_0_stagesList_0_isFlushed;
  wire                DispatchPlugin_logic_pop_0_stagesList_1_isFlushed;
  reg                 DispatchPlugin_logic_pop_0_stagesList_1_LATENCY_0;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_0;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_1;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_2;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_3;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_4;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_5;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_PHYS_RD;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_4;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_5;
  wire                DispatchPlugin_logic_pop_0_stagesList_0_LATENCY_0;
  reg        [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_OFFSET;
  reg        [4:0]    DispatchPlugin_logic_pop_0_stagesList_1_UINT;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID;
  wire       [4:0]    DispatchPlugin_logic_pop_0_stagesList_0_UINT;
  wire                DispatchPlugin_logic_pop_0_stagesList_0_ready;
  wire       [5:0]    DispatchPlugin_logic_pop_0_stagesList_0_OFFSET;
  wire       [31:0]   DispatchPlugin_logic_pop_0_stagesList_0_OH;
  reg        [5:0]    FrontendPlugin_dispatch_PHYS_RS_1_1;
  reg        [5:0]    FrontendPlugin_dispatch_PHYS_RS_0_1;
  reg        [5:0]    FrontendPlugin_dispatch_PHYS_RD_1;
  reg                 FrontendPlugin_dispatch_EU0_SEL_1;
  reg                 FrontendPlugin_dispatch_ALU0_ALU1_SEL_1;
  wire                FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_1;
  reg        [5:0]    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_1;
  wire                FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_1;
  reg        [5:0]    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_1;
  reg                 FrontendPlugin_dispatch_WRITE_RD_1;
  reg        [5:0]    FrontendPlugin_dispatch_PHYS_RS_1_0;
  reg        [5:0]    FrontendPlugin_dispatch_PHYS_RS_0_0;
  reg        [5:0]    FrontendPlugin_dispatch_PHYS_RD_0;
  reg                 FrontendPlugin_dispatch_EU0_SEL_0;
  reg                 FrontendPlugin_dispatch_ALU0_ALU1_SEL_0;
  wire                FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_0;
  wire       [5:0]    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0;
  wire                FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_0;
  wire       [5:0]    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0;
  reg                 FrontendPlugin_dispatch_WRITE_RD_0;
  reg                 FrontendPlugin_dispatch_DispatchPlugin_FENCE_YOUNGER_1;
  reg                 FrontendPlugin_dispatch_DispatchPlugin_FENCE_YOUNGER_0;
  reg                 FrontendPlugin_dispatch_DispatchPlugin_FENCE_OLDER_1;
  reg                 FrontendPlugin_dispatch_DispatchPlugin_FENCE_OLDER_0;
  reg        [1:0]    FrontendPlugin_dispatch_GSHARE_COUNTER_1_0;
  reg        [1:0]    FrontendPlugin_dispatch_GSHARE_COUNTER_1_1;
  reg        [23:0]   FrontendPlugin_dispatch_BRANCH_HISTORY_1;
  reg        [3:0]    FrontendPlugin_dispatch_BRANCH_ID_1;
  reg                 FrontendPlugin_dispatch_BRANCH_SEL_1;
  reg                 _zz_io_writes_1_valid;
  reg        [1:0]    FrontendPlugin_dispatch_GSHARE_COUNTER_0_0;
  reg        [1:0]    FrontendPlugin_dispatch_GSHARE_COUNTER_0_1;
  reg        [23:0]   FrontendPlugin_dispatch_BRANCH_HISTORY_0;
  reg        [3:0]    FrontendPlugin_dispatch_BRANCH_ID_0;
  reg                 FrontendPlugin_dispatch_BRANCH_SEL_0;
  reg                 _zz_io_writes_0_valid;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_isFlushed;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_1_isFlushed;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_isThrown;
  wire                EU0_ExecutionUnitBase_pipeline_execute_1_isFlushed;
  wire                EU0_ExecutionUnitBase_pipeline_execute_2_isFlushed;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E2;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E2;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E2;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_execute_1_PHYS_RD;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_WRITE_RD;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_CsrAccessPlugin_SEL;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_Frontend_MICRO_OP;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_PC;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_VMA;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_VMA;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_VMA;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FLUSH_DATA;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FLUSH_DATA;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FLUSH_DATA;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_I;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_I;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_I;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_XRET;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_XRET;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_XRET;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_ECALL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_ECALL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_ECALL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_EBREAK;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_EBREAK;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_EBREAK;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_HIGH;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_HIGH;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_HIGH;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_CLEAR;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_MASK;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_IMM;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LOAD;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LR;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_PC;
  reg        [4:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_LSU_ID;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_AMO;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SC;
  reg        [0:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_MSB;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SEL;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_REM;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS2_SIGNED;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS1_SIGNED;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS2;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS1;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_completion_SEL_E2;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_execute_2_PHYS_RD;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL;
  wire       [0:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB;
  wire       [4:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_ready;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_isFlushed;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_1_isFlushed;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_isFlushed;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_1_isFlushed;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E1;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E1;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E0;
  reg        [5:0]    ALU1_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  reg        [5:0]    ALU1_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  reg        [3:0]    ALU1_ExecutionUnitBase_pipeline_fetch_1_BRANCH_ID;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_1_PC;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP;
  reg        [1:0]    ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_SEL;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SIGNED;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_LEFT;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SEL;
  reg        [1:0]    ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL;
  reg        [1:0]    ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_SEL;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  reg                 ALU1_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E1;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E0;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_ready;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_WRITE_RD;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire       [1:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL;
  wire       [1:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
  wire       [1:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL;
  wire       [3:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_isFlushed;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_1_isFlushed;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_isFlushed;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_1_isFlushed;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E1;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E1;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E0;
  reg        [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  reg        [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  reg        [3:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_BRANCH_ID;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_1_PC;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP;
  reg        [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_SEL;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SIGNED;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_LEFT;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SEL;
  reg        [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL;
  reg        [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_SEL;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  reg                 ALU0_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E1;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E0;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_ready;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL;
  wire       [3:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
  reg                 FrontendPlugin_dispatch_Prediction_IS_BRANCH_1;
  reg                 FrontendPlugin_dispatch_Prediction_IS_BRANCH_0;
  reg                 FrontendPlugin_serialized_Prediction_IS_BRANCH_1;
  reg                 FrontendPlugin_serialized_Prediction_IS_BRANCH_0;
  wire       [3:0]    FrontendPlugin_serialized_DecoderPredictionPlugin_RAS_PUSH_PTR_1;
  reg                 FrontendPlugin_serialized_RAS_POP_1;
  reg                 DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_2;
  reg                 FrontendPlugin_serialized_RAS_PUSH_1;
  reg        [31:0]   FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_PC_NEXT_1;
  reg                 FrontendPlugin_serialized_BRANCH_EARLY_1_taken;
  reg        [31:0]   FrontendPlugin_serialized_BRANCH_EARLY_1_pc;
  wire                FrontendPlugin_serialized_BRANCH_SEL_1;
  reg                 FrontendPlugin_serialized_CAN_IMPROVE_1;
  reg                 FrontendPlugin_serialized_Frontend_DECODED_MASK_1;
  wire                FrontendPlugin_serialized_NEED_CORRECTION_1;
  wire                FrontendPlugin_serialized_MISSMATCH_1;
  wire                FrontendPlugin_serialized_MISSMATCH_HISTORY_1;
  reg                 FrontendPlugin_serialized_BAD_RET_PC_1;
  wire                FrontendPlugin_serialized_MISSMATCH_PC_1;
  reg                 FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_1;
  reg                 FrontendPlugin_serialized_IS_ANY_1;
  reg        [31:0]   FrontendPlugin_serialized_PC_INC_1;
  reg                 FrontendPlugin_serialized_BRANCHED_PREDICTION_1;
  wire       [31:0]   FrontendPlugin_serialized_PC_PREDICTION_1;
  reg                 FrontendPlugin_serialized_IS_JALR_1;
  reg        [31:0]   FrontendPlugin_serialized_PC_TARGET_PRE_RAS_1;
  reg        [31:0]   FrontendPlugin_serialized_PC_TARGET_1;
  wire                FrontendPlugin_decoded_BRANCHED_PREDICTION_1;
  wire                FrontendPlugin_decoded_CAN_IMPROVE_1;
  wire       [31:0]   FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_1;
  wire                FrontendPlugin_decoded_BAD_RET_PC_1;
  wire       [31:0]   FrontendPlugin_decoded_PC_TARGET_PRE_RAS_1;
  wire       [31:0]   FrontendPlugin_decoded_PC_INC_1;
  wire       [1:0]    FrontendPlugin_decoded_Prediction_CONDITIONAL_TAKE_IT_1;
  wire                FrontendPlugin_decoded_CONDITIONAL_PREDICTION_1;
  wire       [0:0]    FrontendPlugin_decoded_LAST_SLICE_1;
  wire                FrontendPlugin_decoded_RAS_POP_1;
  wire                FrontendPlugin_decoded_RAS_PUSH_1;
  wire       [31:0]   FrontendPlugin_decoded_OFFSET_1;
  wire                FrontendPlugin_decoded_IS_ANY_1;
  wire                FrontendPlugin_decoded_Prediction_IS_BRANCH_1;
  wire                FrontendPlugin_decoded_IS_JALR_1;
  wire                FrontendPlugin_decoded_IS_JAL_1;
  wire       [3:0]    FrontendPlugin_serialized_DecoderPredictionPlugin_RAS_PUSH_PTR_0;
  reg                 FrontendPlugin_serialized_RAS_POP_0;
  reg                 DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_1;
  reg                 FrontendPlugin_serialized_RAS_PUSH_0;
  reg        [31:0]   FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  reg                 FrontendPlugin_serialized_BRANCH_EARLY_0_taken;
  reg        [31:0]   FrontendPlugin_serialized_BRANCH_EARLY_0_pc;
  wire                FrontendPlugin_serialized_BRANCH_SEL_0;
  reg                 FrontendPlugin_serialized_CAN_IMPROVE_0;
  reg                 FrontendPlugin_serialized_Frontend_DECODED_MASK_0;
  wire                FrontendPlugin_serialized_NEED_CORRECTION_0;
  wire                FrontendPlugin_serialized_MISSMATCH_0;
  wire                FrontendPlugin_serialized_MISSMATCH_HISTORY_0;
  reg                 FrontendPlugin_serialized_BAD_RET_PC_0;
  wire                FrontendPlugin_serialized_MISSMATCH_PC_0;
  reg                 FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0;
  reg                 FrontendPlugin_serialized_IS_ANY_0;
  reg        [31:0]   FrontendPlugin_serialized_PC_INC_0;
  reg                 FrontendPlugin_serialized_BRANCHED_PREDICTION_0;
  wire       [31:0]   FrontendPlugin_serialized_PC_PREDICTION_0;
  reg                 FrontendPlugin_serialized_IS_JALR_0;
  reg        [31:0]   FrontendPlugin_serialized_PC_TARGET_PRE_RAS_0;
  reg        [31:0]   FrontendPlugin_serialized_PC_TARGET_0;
  wire                FrontendPlugin_decoded_BRANCHED_PREDICTION_0;
  wire                FrontendPlugin_decoded_CAN_IMPROVE_0;
  wire       [31:0]   FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  wire                FrontendPlugin_decoded_BAD_RET_PC_0;
  wire       [31:0]   FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0;
  wire       [31:0]   FrontendPlugin_decoded_PC_INC_0;
  wire       [1:0]    FrontendPlugin_decoded_Prediction_CONDITIONAL_TAKE_IT_0;
  wire                FrontendPlugin_decoded_CONDITIONAL_PREDICTION_0;
  wire       [0:0]    FrontendPlugin_decoded_LAST_SLICE_0;
  wire                FrontendPlugin_decoded_RAS_POP_0;
  wire                FrontendPlugin_decoded_RAS_PUSH_0;
  wire       [31:0]   FrontendPlugin_decoded_OFFSET_0;
  wire                FrontendPlugin_decoded_IS_ANY_0;
  wire                FrontendPlugin_decoded_Prediction_IS_BRANCH_0;
  wire                FrontendPlugin_decoded_IS_JALR_0;
  reg        [31:0]   FrontendPlugin_dispatch_Frontend_MICRO_OP_1;
  wire                FrontendPlugin_dispatch_LATENCY_0_1;
  reg        [31:0]   FrontendPlugin_dispatch_Frontend_MICRO_OP_0;
  wire                FrontendPlugin_dispatch_LATENCY_0_0;
  wire       [11:0]   FrontendPlugin_allocated_OP_ID /* verilator public */ ;
  reg        [11:0]   FrontendPlugin_decoded_OP_ID /* verilator public */ ;
  wire       [3:0]    FrontendPlugin_allocated_DecoderPredictionPlugin_RAS_PUSH_PTR_1;
  wire       [3:0]    FrontendPlugin_allocated_DecoderPredictionPlugin_RAS_PUSH_PTR_0;
  wire       [31:0]   FrontendPlugin_allocated_Frontend_MICRO_OP_1;
  wire       [31:0]   FrontendPlugin_allocated_Frontend_MICRO_OP_0;
  wire                FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_1;
  wire                FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_1;
  wire                FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1;
  reg        [31:0]   FrontendPlugin_serialized_Frontend_MICRO_OP_1;
  wire                FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1;
  wire                FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0;
  wire                FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0;
  wire                FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0;
  reg        [31:0]   FrontendPlugin_serialized_Frontend_MICRO_OP_0;
  wire                FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0;
  wire       [31:0]   FrontendPlugin_decoded_Frontend_INSTRUCTION_ALIGNED_1;
  wire       [31:0]   FrontendPlugin_decoded_Frontend_INSTRUCTION_ALIGNED_0;
  wire       [31:0]   FrontendPlugin_decoded_PC_1 /* verilator public */ ;
  wire       [31:0]   FrontendPlugin_decoded_PC_0 /* verilator public */ ;
  wire                FrontendPlugin_decoded_Frontend_FETCH_FAULT_PAGE_1;
  wire                FrontendPlugin_decoded_Frontend_FETCH_FAULT_PAGE_0;
  wire                FrontendPlugin_decoded_isFlushed;
  wire       [4:0]    FrontendPlugin_decoded_ARCH_RS_1_1;
  wire       [4:0]    FrontendPlugin_decoded_ARCH_RS_0_1;
  wire       [4:0]    FrontendPlugin_decoded_ARCH_RD_1;
  wire       [31:0]   FrontendPlugin_decoded_Frontend_MICRO_OP_1;
  wire                FrontendPlugin_decoded_Frontend_DECODED_MASK_1 /* verilator public */ ;
  wire                FrontendPlugin_decoded_Frontend_FETCH_FAULT_1;
  wire                FrontendPlugin_decoded_Frontend_MASK_ALIGNED_1;
  wire                FrontendPlugin_decoded_TRAP_1;
  wire                FrontendPlugin_decoded_SQ_ALLOC_1;
  wire                FrontendPlugin_decoded_LQ_ALLOC_1;
  wire                FrontendPlugin_decoded_EU0_SEL_1;
  wire                FrontendPlugin_decoded_ALU0_ALU1_SEL_1;
  wire                FrontendPlugin_decoded_WRITE_RD_1;
  wire                FrontendPlugin_decoded_READ_RS_1_1;
  wire                FrontendPlugin_decoded_READ_RS_0_1;
  wire                FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_1;
  wire                FrontendPlugin_decoded_LEGAL_1;
  wire       [31:0]   FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 /* verilator public */ ;
  wire       [4:0]    FrontendPlugin_decoded_ARCH_RS_1_0;
  wire       [4:0]    FrontendPlugin_decoded_ARCH_RS_0_0;
  wire       [4:0]    FrontendPlugin_decoded_ARCH_RD_0;
  wire       [31:0]   FrontendPlugin_decoded_Frontend_MICRO_OP_0;
  wire                FrontendPlugin_decoded_Frontend_DECODED_MASK_0 /* verilator public */ ;
  wire                FrontendPlugin_decoded_Frontend_FETCH_FAULT_0;
  wire                FrontendPlugin_decoded_Frontend_MASK_ALIGNED_0;
  wire                FrontendPlugin_decoded_TRAP_0;
  wire                FrontendPlugin_decoded_SQ_ALLOC_0;
  wire                FrontendPlugin_decoded_LQ_ALLOC_0;
  wire                FrontendPlugin_decoded_EU0_SEL_0;
  wire                FrontendPlugin_decoded_ALU0_ALU1_SEL_0;
  wire                FrontendPlugin_decoded_WRITE_RD_0;
  wire                FrontendPlugin_decoded_READ_RS_1_0;
  wire                FrontendPlugin_decoded_READ_RS_0_0;
  wire                FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_0;
  wire                FrontendPlugin_decoded_LEGAL_0;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_CLEAR;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_IMM;
  reg                 _zz_9;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_isFlushed;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_isThrown;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_isFlushed;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_isThrown;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_isFlushed;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_isThrown;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_isFlushed;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_isFlushed;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_isFlushed;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH_PC;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH_PC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_SP_FP_ADDRESS;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_SP_FP_ADDRESS;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION_COUNTER;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION_COUNTER;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_AMO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_AMO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_SC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_SC;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_DELTA;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_DELTA;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_VALID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_VALID;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SCORE;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SCORE;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_MMU_TRANSLATED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LR;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LR;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_2_SQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_1_PHYS_RD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_WRITE_RD;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_1_ROB_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_UNSIGNED;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_1_SIZE;
  reg                 FetchPlugin_stages_1_MMU_ACCESS_FAULT;
  reg                 FetchPlugin_stages_1_MMU_PAGE_FAULT;
  reg                 FetchPlugin_stages_1_MMU_ALLOW_WRITE;
  reg                 FetchPlugin_stages_1_MMU_ALLOW_READ;
  reg                 FetchPlugin_stages_1_MMU_ALLOW_EXECUTE;
  reg                 FetchPlugin_stages_1_MMU_REDO;
  reg        [31:0]   FetchPlugin_stages_1_MMU_TRANSLATED;
  wire                FetchPlugin_stages_1_MMU_IO;
  reg        [1:0]    FetchPlugin_stages_1_MMU_L1_HITS;
  reg        [1:0]    FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_pageFault;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_accessFault;
  wire       [4:0]    FetchPlugin_stages_1_MMU_L1_ENTRIES_0_virtualAddress;
  wire       [9:0]    FetchPlugin_stages_1_MMU_L1_ENTRIES_0_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowRead;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowUser;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_pageFault;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_accessFault;
  wire       [4:0]    FetchPlugin_stages_1_MMU_L1_ENTRIES_1_virtualAddress;
  wire       [9:0]    FetchPlugin_stages_1_MMU_L1_ENTRIES_1_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowRead;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowUser;
  reg        [3:0]    FetchPlugin_stages_1_MMU_L0_HITS;
  reg        [3:0]    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_pageFault;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_accessFault;
  wire       [14:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_0_virtualAddress;
  wire       [19:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_0_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowRead;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowUser;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_pageFault;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_accessFault;
  wire       [14:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_1_virtualAddress;
  wire       [19:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_1_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowRead;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowUser;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_pageFault;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_accessFault;
  wire       [14:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_2_virtualAddress;
  wire       [19:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_2_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowRead;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowUser;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_pageFault;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_accessFault;
  wire       [14:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_3_virtualAddress;
  wire       [19:0]   FetchPlugin_stages_1_MMU_L0_ENTRIES_3_physicalAddress;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowRead;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowWrite;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowExecute;
  wire                FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowUser;
  wire                FetchPlugin_stages_1_isRemoved;
  wire                FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded;
  wire                FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_0;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_1;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_2;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_3;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_4;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_5;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_OH;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_MMU_BYPASS_TRANSLATION;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_WRITE;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_EXECUTE;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_accessFault;
  reg        [4:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_virtualAddress;
  reg        [9:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_accessFault;
  reg        [4:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_virtualAddress;
  reg        [9:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowUser;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS_PRE_VALID;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_HITS_PRE_VALID;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_accessFault;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_virtualAddress;
  wire       [9:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_accessFault;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_virtualAddress;
  wire       [9:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_accessFault;
  reg        [14:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_virtualAddress;
  reg        [19:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_accessFault;
  reg        [14:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_virtualAddress;
  reg        [19:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_accessFault;
  reg        [14:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_virtualAddress;
  reg        [19:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowUser;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_pageFault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_accessFault;
  reg        [14:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_virtualAddress;
  reg        [19:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_physicalAddress;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowRead;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowWrite;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowExecute;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowUser;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_accessFault;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_virtualAddress;
  wire       [19:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_accessFault;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_virtualAddress;
  wire       [19:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_accessFault;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_virtualAddress;
  wire       [19:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_pageFault;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_accessFault;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_virtualAddress;
  wire       [19:0]   Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_physicalAddress;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowRead;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowWrite;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowExecute;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowUser;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_isRemoved;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_isRemoved;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL_overloaded;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_1_PC_TRUE;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_1_PC;
  reg        [3:0]    ALU1_ExecutionUnitBase_pipeline_execute_1_BRANCH_ID;
  reg                 _zz_io_writes_1_valid_1;
  reg                 ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_1_ready;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED;
  reg        [1:0]    ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_1_PC_TARGET;
  reg        [5:0]    ALU1_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
  reg                 ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BAD_EARLY_TARGET;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSPREDICTED;
  reg                 ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND;
  reg                 ALU1_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_taken;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_pc;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BAD_EARLY_TARGET;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_1_PC_TRUE;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_1_PC;
  reg        [3:0]    ALU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_ID;
  reg                 _zz_io_writes_0_valid_1;
  reg                 ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_1_ready;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED;
  reg        [1:0]    ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET;
  reg        [5:0]    ALU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
  reg                 ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BAD_EARLY_TARGET;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSPREDICTED;
  reg                 ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND;
  reg                 ALU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_taken;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_pc;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BAD_EARLY_TARGET;
  reg                 _zz_FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH_PC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_SP_FP_ADDRESS;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION_COUNTER;
  reg                 _zz_io_writes_2_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_AMO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_SC;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ROB;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_DELTA;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_VALID;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE;
  reg                 _zz_io_writes_2_valid_1;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_MMU_TRANSLATED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LR;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_WRITE_RD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_IS_IO;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_resulting;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_resulting;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_WAIT_FEED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_ready;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_3_CTRL;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_valid;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_data;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_fault;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlot;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlotAny;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_ADDRESS_PRE_TRANSLATION;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_3_PHYS_RD;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ID;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_valid;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_data;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_fault;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_redo;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlot;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_valid;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_data;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_fault;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlot;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_valid;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_data;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_fault;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlot;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_TRAP_SPECULATION;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_2_CTRL;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_WRITE;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_PAGE_FAULT;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_MISS_ALIGNED;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_WRITE_FAILURE;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_2_PHYS_RD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_ACCESS_FAULT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_READ;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_WRITE_RD;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_2_LQ_ID;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_MMU_REDO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_IS_IO;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_ready;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_HIT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_UNSIGNED;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_valid;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_fault;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlot;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlotAny;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ID;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_RESCHEDULE;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ROB;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_NO_YOUNGER;
  reg        [15:0]   Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER;
  reg        [15:0]   Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS;
  reg        [4:0]    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_BYPASS_SUCCESS;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_2_SIZE;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_TRANSLATED;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_overloaded;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED_overloaded;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED;
  reg                 _zz_io_writes_1_valid_2;
  reg                 _zz_10;
  reg                 _zz_11;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID;
  reg                 _zz_io_writes_1_valid_3;
  reg                 _zz_12;
  reg                 _zz_13;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_ready;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_OH;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_ID;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_HIT;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_NO_OLDER;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK;
  reg        [4:0]    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID;
  reg        [4:0]    Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_TRANSLATED_AS_IO;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_IS_IO;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_POST_TRANSLATION;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION;
  reg                 _zz_io_writes_2_valid_2;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH_PC;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SQID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SQID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SQID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_FEEDED;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SQID;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_stages_0_feed_SQ_PTR_FREE;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_stages_0_SQCHECK_END_ID;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_stages_0_LQCHECK_START_ID;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD_agu;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD_agu;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_agu;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_SP_FP_ADDRESS;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION_COUNTER;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_SC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_AMO;
  reg        [2:0]    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SCORE;
  reg        [3:0]    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID;
  reg        [4:0]    Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_LR;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_UNSIGNED;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_store;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_load;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_store;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_load;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_stages_0_SIZE;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_0_SIZE_store;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_stages_0_SIZE_load;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_store;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_load;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_store;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_load;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s1_ready;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_isRemoved;
  reg                 _zz_Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_ready;
  wire       [6:0]    Lsu2Plugin_logic_sharedPip_stages_0_SQ_ROB_FULL;
  wire       [6:0]    Lsu2Plugin_logic_sharedPip_stages_0_LQ_ROB_FULL;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ;
  reg        [3:0]    Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID;
  reg        [3:0]    Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID;
  reg                 Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s1_LQ_HIT;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s1_SQ_HIT;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_LQ_OLDER_THAN_SQ;
  reg        [6:0]    Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ROB_FULL;
  reg        [6:0]    Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ROB_FULL;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_ready;
  wire       [6:0]    Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ROB_FULL;
  wire       [6:0]    Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ROB_FULL;
  wire       [3:0]    Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID;
  wire       [3:0]    Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH;
  reg        [5:0]    FrontendPlugin_dispatch_ROB_ID /* verilator public */ ;
  reg        [4:0]    Lsu2Plugin_logic_allocation_stores_alloc_2;
  reg                 _zz_io_writes_1_valid_4;
  reg                 _zz_io_writes_1_valid_5;
  reg                 _zz_io_writes_1_valid_6;
  reg        [4:0]    Lsu2Plugin_logic_allocation_loads_alloc_2;
  reg                 _zz_14;
  reg        [4:0]    FrontendPlugin_dispatch_ARCH_RS_0_1;
  reg                 _zz_io_writes_1_valid_7;
  reg                 _zz_io_writes_1_valid_8;
  wire       [3:0]    FrontendPlugin_dispatch_SQ_ID_1;
  wire       [3:0]    FrontendPlugin_dispatch_LQ_ID_1;
  reg        [4:0]    Lsu2Plugin_logic_allocation_stores_alloc_1;
  reg                 _zz_io_writes_0_valid_2;
  reg                 _zz_io_writes_0_valid_3;
  reg                 _zz_io_writes_0_valid_4;
  reg        [4:0]    Lsu2Plugin_logic_allocation_loads_alloc_1;
  reg                 _zz_15;
  reg        [4:0]    FrontendPlugin_dispatch_ARCH_RS_0_0;
  reg                 _zz_io_writes_0_valid_5;
  reg                 _zz_io_writes_0_valid_6;
  reg                 FrontendPlugin_dispatch_ready;
  wire       [3:0]    FrontendPlugin_dispatch_SQ_ID_0;
  wire       [3:0]    FrontendPlugin_dispatch_LQ_ID_0;
  reg                 FrontendPlugin_dispatch_SQ_ALLOC_1;
  reg                 FrontendPlugin_dispatch_SQ_ALLOC_0;
  reg                 FrontendPlugin_dispatch_LQ_ALLOC_1;
  reg                 FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1 /* verilator public */ ;
  reg                 FrontendPlugin_dispatch_LQ_ALLOC_0;
  reg                 FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 /* verilator public */ ;
  reg        [4:0]    FrontendPlugin_dispatch_LSU_ID_1;
  reg        [4:0]    FrontendPlugin_dispatch_LSU_ID_0;
  reg        [4:0]    Lsu2Plugin_logic_sq_onCommit_commitComb_2;
  reg        [4:0]    Lsu2Plugin_logic_sq_onCommit_commitComb_1;
  reg                 _zz_when_MultiportRam_l362;
  reg                 _zz_when_MultiportRam_l362_1;
  reg        [4:0]    Lsu2Plugin_logic_lq_onCommit_free_2;
  reg        [14:0]   Lsu2Plugin_logic_lq_onCommit_priority_2;
  reg        [4:0]    Lsu2Plugin_logic_lq_onCommit_free_1;
  reg        [14:0]   Lsu2Plugin_logic_lq_onCommit_priority_1;
  wire       [31:0]   FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 /* verilator public */ ;
  wire                FrontendPlugin_decoded_IS_JAL_0;
  wire       [23:0]   FrontendPlugin_allocated_BRANCH_HISTORY_1 /* verilator public */ ;
  wire       [23:0]   FrontendPlugin_allocated_BRANCH_HISTORY_0 /* verilator public */ ;
  reg        [23:0]   HistoryPlugin_logic_update_pushes_2_stateNext_2;
  reg        [23:0]   HistoryPlugin_logic_update_pushes_2_stateNext_1;
  reg        [23:0]   HistoryPlugin_logic_update_pushes_0_stateNext_1;
  reg        [23:0]   HistoryPlugin_logic_onCommit_valueNext_2;
  reg        [23:0]   HistoryPlugin_logic_onCommit_valueNext_1;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RS_1_1;
  wire                FrontendPlugin_allocated_READ_RS_1_1;
  wire       [4:0]    FrontendPlugin_allocated_ARCH_RS_1_1;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RS_0_1;
  wire                FrontendPlugin_allocated_READ_RS_0_1;
  wire       [4:0]    FrontendPlugin_allocated_ARCH_RS_0_1;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RD_FREE_1;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RS_1_0;
  wire                FrontendPlugin_allocated_READ_RS_1_0;
  wire       [4:0]    FrontendPlugin_allocated_ARCH_RS_1_0;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RS_0_0;
  wire                FrontendPlugin_allocated_READ_RS_0_0;
  wire       [4:0]    FrontendPlugin_allocated_ARCH_RS_0_0;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RD_FREE_0;
  wire       [4:0]    FrontendPlugin_allocated_ARCH_RD_1;
  wire       [4:0]    FrontendPlugin_allocated_ARCH_RD_0;
  wire       [3:0]    ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TARGET;
  (* keep , syn_keep *) wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TRUE /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_PC;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
  wire       [1:0]    ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SHIFT_RESULT;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SIGNED;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SEL;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_RESULT;
  wire       [1:0]    ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL;
  wire       [1:0]    ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_SEL;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
  wire       [1:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
  wire       [0:0]    ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC1_CTRL;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_ready;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_2_Frontend_MICRO_OP;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_2_PC;
  reg        [5:0]    EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LOAD;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LR;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_PC;
  wire       [4:0]    EU0_ExecutionUnitBase_pipeline_execute_0_LSU_ID;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_AMO;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SC;
  wire       [0:0]    EU0_ExecutionUnitBase_pipeline_execute_0_ROB_MSB;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_isRemoved;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_DIV_RESULT;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_DIV_REVERT_RESULT;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_REM;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_ready;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_0_ready;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_DIV_REVERT_RESULT;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_HIGH;
  wire       [65:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0;
  reg        [4:0]    EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_0_adders_1;
  reg        [62:0]   EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_0_adders_0;
  wire       [4:0]    EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1;
  wire       [62:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0;
  reg        [46:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_2;
  reg        [46:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_1;
  reg        [29:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_3;
  reg        [33:0]   EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_0;
  (* keep , syn_keep *) wire       [29:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [46:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [46:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [33:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [32:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [32:0]   EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1 /* synthesis syn_keep = 1 */ ;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_SIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
  wire       [0:0]    EU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  wire       [3:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TARGET;
  (* keep , syn_keep *) wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_PC;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SHIFT_RESULT;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SIGNED;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SEL;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_RESULT;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_SEL;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
  wire       [1:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
  wire       [0:0]    ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC1_CTRL;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  wire       [31:0]   FrontendPlugin_allocated_PC_1;
  wire       [31:0]   FrontendPlugin_allocated_PC_0;
  reg                 CommitPlugin_logic_commit_continue_2;
  reg                 CommitPlugin_logic_commit_continue_1;
  wire       [0:0]    FrontendPlugin_allocated_ROB_MSB_1;
  wire       [0:0]    FrontendPlugin_allocated_ROB_MSB_0;
  wire       [1:0]    FrontendPlugin_decompressed_GSHARE_COUNTER_1_0;
  wire       [1:0]    FrontendPlugin_decompressed_GSHARE_COUNTER_1_1;
  wire       [1:0]    FrontendPlugin_decompressed_Prediction_CONDITIONAL_TAKE_IT_1;
  wire       [1:0]    FrontendPlugin_decompressed_GSHARE_COUNTER_0_0;
  wire       [1:0]    FrontendPlugin_decompressed_GSHARE_COUNTER_0_1;
  wire       [1:0]    FrontendPlugin_decompressed_Prediction_CONDITIONAL_TAKE_IT_0;
  reg        [12:0]   FetchPlugin_stages_1_GSharePlugin_logic_HASH;
  reg                 FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_valid;
  reg        [12:0]   FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_address;
  reg        [1:0]    FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_data_0;
  reg        [1:0]    FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_data_1;
  wire                FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_valid;
  wire       [12:0]   FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_data_0;
  wire       [1:0]    FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_data_1;
  wire       [23:0]   FetchPlugin_stages_0_BRANCH_HISTORY;
  wire       [12:0]   FetchPlugin_stages_0_GSharePlugin_logic_HASH;
  reg                 _zz_when_MultiportRam_l328;
  wire                FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALUE;
  wire       [0:0]    FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_SLICE;
  wire                FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALID;
  wire       [31:0]   FetchPlugin_stages_1_Prediction_WORD_BRANCH_PC_NEXT;
  wire       [0:0]    FetchPlugin_stages_1_Prediction_WORD_BRANCH_SLICE;
  wire                FetchPlugin_stages_1_Prediction_WORD_BRANCH_VALID;
  (* keep , syn_keep *) reg        [1:0]    FetchPlugin_stages_1_GSHARE_COUNTER_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    FetchPlugin_stages_1_GSHARE_COUNTER_1 /* synthesis syn_keep = 1 */ ;
  wire                FetchPlugin_stages_1_BtbPlugin_logic_HIT;
  (* keep , syn_keep *) wire       [15:0]   FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [0:0]    FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_slice /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_pcTarget /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_isBranch /* synthesis syn_keep = 1 */ ;
  reg                 _zz_16;
  reg                 _zz_17;
  wire       [5:0]    FrontendPlugin_allocated_ROB_ID /* verilator public */ ;
  reg                 _zz_io_writes_1_valid_9;
  wire                FrontendPlugin_allocated_BRANCH_EARLY_1_taken;
  wire       [31:0]   FrontendPlugin_allocated_BRANCH_EARLY_1_pc;
  reg        [4:0]    BranchContextPlugin_logic_alloc_allocNext_2;
  wire                FrontendPlugin_allocated_BRANCH_SEL_1;
  wire       [3:0]    FrontendPlugin_allocated_BRANCH_ID_1;
  reg                 _zz_io_writes_0_valid_7;
  wire                FrontendPlugin_allocated_BRANCH_EARLY_0_taken;
  wire       [31:0]   FrontendPlugin_allocated_BRANCH_EARLY_0_pc;
  reg        [4:0]    BranchContextPlugin_logic_alloc_allocNext_1;
  wire                FrontendPlugin_allocated_BRANCH_SEL_0;
  wire       [3:0]    FrontendPlugin_allocated_BRANCH_ID_0;
  wire                FrontendPlugin_serialized_isFlushed;
  reg                 FrontendPlugin_serialized_ready;
  wire                FrontendPlugin_serialized_isForked;
  wire                FrontendPlugin_serialized_Frontend_DISPATCH_MASK_1_overloaded;
  wire                FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0_overloaded;
  wire                FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_1;
  wire                FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0;
  wire                FrontendPlugin_serialized_Frontend_DISPATCH_MASK_1;
  wire                FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RD_1;
  wire                FrontendPlugin_allocated_WRITE_RD_1;
  wire                FrontendPlugin_allocated_Frontend_DISPATCH_MASK_1;
  reg        [5:0]    FrontendPlugin_allocated_PHYS_RD_0;
  wire                FrontendPlugin_allocated_WRITE_RD_0;
  wire                FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0;
  wire                FrontendPlugin_decompressed_Frontend_INSTRUCTION_ILLEGAL_1;
  wire       [31:0]   FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_1;
  wire       [31:0]   FrontendPlugin_decompressed_Frontend_INSTRUCTION_DECOMPRESSED_1;
  wire                FrontendPlugin_decompressed_Frontend_INSTRUCTION_ILLEGAL_0;
  wire       [31:0]   FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_0;
  wire       [31:0]   FrontendPlugin_decompressed_Frontend_INSTRUCTION_DECOMPRESSED_0;
  wire                FrontendPlugin_aligned_isFlushed;
  reg        [31:0]   AlignerPlugin_setup_s2m_Fetch_FETCH_PC_INC;
  wire                AlignerPlugin_setup_s2m_isFlushed;
  reg                 AlignerPlugin_setup_s2m_ready;
  wire                FrontendPlugin_aligned_ready;
  reg                 FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_1;
  reg                 FrontendPlugin_aligned_Frontend_FETCH_FAULT_1;
  reg        [11:0]   FrontendPlugin_aligned_FETCH_ID_1;
  reg        [1:0]    FrontendPlugin_aligned_GSHARE_COUNTER_1_0;
  reg        [1:0]    FrontendPlugin_aligned_GSHARE_COUNTER_1_1;
  reg                 FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALUE_1;
  reg        [0:0]    FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_SLICE_1;
  reg                 FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALID_1;
  reg        [23:0]   FrontendPlugin_aligned_BRANCH_HISTORY_1;
  reg        [31:0]   FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_1;
  reg                 FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1;
  wire       [31:0]   FrontendPlugin_aligned_PC_1;
  wire                FrontendPlugin_aligned_Frontend_MASK_ALIGNED_1;
  wire       [31:0]   FrontendPlugin_aligned_Frontend_INSTRUCTION_ALIGNED_1;
  reg        [3:0]    AlignerPlugin_logic_slices_remains_2;
  reg        [3:0]    AlignerPlugin_logic_slices_carry_2;
  reg        [3:0]    AlignerPlugin_logic_slices_used_2;
  reg                 AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE;
  reg                 AlignerPlugin_setup_s2m_Fetch_WORD_FAULT;
  reg                 FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0;
  reg                 FrontendPlugin_aligned_Frontend_FETCH_FAULT_0;
  reg        [11:0]   AlignerPlugin_setup_s2m_FETCH_ID;
  reg        [11:0]   FrontendPlugin_aligned_FETCH_ID_0;
  reg        [31:0]   AlignerPlugin_setup_s2m_Fetch_FETCH_PC;
  reg        [1:0]    AlignerPlugin_setup_s2m_GSHARE_COUNTER_0;
  reg        [1:0]    AlignerPlugin_setup_s2m_GSHARE_COUNTER_1;
  reg        [1:0]    FrontendPlugin_aligned_GSHARE_COUNTER_0_0;
  reg        [1:0]    FrontendPlugin_aligned_GSHARE_COUNTER_0_1;
  reg                 AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE;
  reg                 FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALUE_0;
  reg        [0:0]    AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_SLICE;
  reg        [0:0]    FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_SLICE_0;
  reg                 AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID;
  reg                 FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALID_0;
  reg        [23:0]   AlignerPlugin_setup_s2m_BRANCH_HISTORY;
  reg        [23:0]   FrontendPlugin_aligned_BRANCH_HISTORY_0;
  reg        [31:0]   AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT;
  reg        [31:0]   FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  reg                 FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0;
  wire       [31:0]   FrontendPlugin_aligned_PC_0;
  wire                FrontendPlugin_aligned_Frontend_MASK_ALIGNED_0;
  wire       [31:0]   FrontendPlugin_aligned_Frontend_INSTRUCTION_ALIGNED_0;
  reg        [3:0]    AlignerPlugin_logic_slices_remains_1;
  reg        [3:0]    AlignerPlugin_logic_slices_carry_1;
  reg        [3:0]    AlignerPlugin_logic_slices_used_1;
  reg        [1:0]    AlignerPlugin_setup_s2m_MASK_FRONT;
  reg        [63:0]   AlignerPlugin_setup_s2m_Fetch_WORD;
  reg                 AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID;
  reg        [0:0]    AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_SLICE;
  reg        [1:0]    AlignerPlugin_setup_s2m_MASK_BACK;
  wire       [1:0]    FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT;
  wire                AlignerPlugin_setup_s2m_isFlushingRoot;
  reg        [23:0]   FetchPlugin_stages_2_BRANCH_HISTORY;
  reg                 FetchPlugin_stages_2_MMU_IO;
  reg        [31:0]   FetchPlugin_stages_2_MMU_TRANSLATED;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HIT;
  reg                 FetchPlugin_stages_2_MMU_REDO;
  wire                FetchPlugin_stages_2_ready;
  reg                 _zz_FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552;
  reg                 _zz_FetchPlugin_stages_2_isFlushingRoot;
  reg                 FetchPlugin_stages_2_MMU_ALLOW_EXECUTE;
  reg                 FetchPlugin_stages_2_MMU_PAGE_FAULT;
  reg                 FetchPlugin_stages_2_MMU_ACCESS_FAULT;
  wire                FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_error;
  reg        [19:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_address;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_1_loaded;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_1_error;
  reg        [19:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_1_address;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_2_loaded;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_2_error;
  reg        [19:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_2_address;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_3_loaded;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_3_error;
  reg        [19:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_3_address;
  wire                FetchPlugin_stages_2_Fetch_WORD_FAULT;
  reg        [31:0]   FetchPlugin_stages_2_Fetch_FETCH_PC;
  reg        [0:0]    FetchPlugin_stages_2_FetchCachePlugin_logic_PLRU_0;
  reg        [1:0]    FetchPlugin_stages_2_FetchCachePlugin_logic_PLRU_1;
  wire                FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HIT;
  wire       [0:0]    FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0;
  wire       [1:0]    FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_1;
  wire                FetchPlugin_stages_1_MMU_BYPASS_TRANSLATION;
  wire                FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_0;
  wire                FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_1;
  wire                FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_2;
  wire                FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_3;
  wire       [5:0]    FetchPlugin_stages_1_MMU_WAYS_OH;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_0;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_1;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_2;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_3;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_4;
  wire       [31:0]   FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_5;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_error;
  reg        [19:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_loaded;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_error;
  reg        [19:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_loaded;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_error;
  reg        [19:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_loaded;
  reg                 FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_error;
  reg        [19:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address;
  reg        [63:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_0;
  reg        [63:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_1;
  reg        [63:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_2;
  reg        [63:0]   FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_3;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_0;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_1;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_2;
  reg                 FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_3;
  wire       [63:0]   FetchPlugin_stages_2_Fetch_WORD;
  reg        [31:0]   FetchPlugin_stages_1_Fetch_FETCH_PC;
  wire       [63:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_0;
  wire       [63:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_1;
  wire       [63:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_2;
  wire       [63:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_3;
  wire       [31:0]   FetchPlugin_stages_0_Fetch_FETCH_PC;
  reg                 FetchPlugin_stages_0_ready;
  reg                 _zz_18;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_error;
  wire       [19:0]   FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_address;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_1_loaded;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_1_error;
  wire       [19:0]   FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_1_address;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_2_loaded;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_2_error;
  wire       [19:0]   FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_2_address;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_3_loaded;
  wire                FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_3_error;
  wire       [19:0]   FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_3_address;
  reg                 _zz_when_MultiportRam_l328_1;
  reg                 _zz_when_MultiportRam_l328_2;
  reg                 _zz_when_MultiportRam_l328_3;
  wire       [63:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_0;
  wire       [63:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_1;
  wire       [63:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_2;
  wire       [63:0]   FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_3;
  reg                 _zz_when_MultiportRam_l328_4;
  reg        [31:0]   PcPlugin_logic_jump_target_1;
  wire                FetchPlugin_stages_1_isFlushed;
  wire                FetchPlugin_stages_1_ready;
  reg        [11:0]   FetchPlugin_stages_1_FETCH_ID /* verilator public */ ;
  wire       [11:0]   FrontendPlugin_allocated_FETCH_ID_1 /* verilator public */ ;
  wire       [11:0]   FrontendPlugin_decoded_FETCH_ID_1 /* verilator public */ ;
  reg                 FrontendPlugin_allocated_ready;
  reg                 FrontendPlugin_decoded_ready;
  wire       [11:0]   FrontendPlugin_allocated_FETCH_ID_0 /* verilator public */ ;
  wire       [11:0]   FrontendPlugin_decoded_FETCH_ID_0 /* verilator public */ ;
  reg                 MmuPlugin_setup_cacheLoad_cmd_valid;
  wire                MmuPlugin_setup_cacheLoad_cmd_ready;
  wire       [31:0]   MmuPlugin_setup_cacheLoad_cmd_payload_virtual;
  wire       [1:0]    MmuPlugin_setup_cacheLoad_cmd_payload_size;
  wire                MmuPlugin_setup_cacheLoad_cmd_payload_redoOnDataHazard;
  wire                MmuPlugin_setup_cacheLoad_cmd_payload_unlocked;
  wire                MmuPlugin_setup_cacheLoad_cmd_payload_unique;
  wire       [31:0]   MmuPlugin_setup_cacheLoad_translated_physical;
  wire                MmuPlugin_setup_cacheLoad_translated_abord;
  wire       [2:0]    MmuPlugin_setup_cacheLoad_cancels;
  wire                MmuPlugin_setup_cacheLoad_rsp_valid;
  wire       [31:0]   MmuPlugin_setup_cacheLoad_rsp_payload_data;
  wire                MmuPlugin_setup_cacheLoad_rsp_payload_fault;
  wire                MmuPlugin_setup_cacheLoad_rsp_payload_redo;
  wire       [1:0]    MmuPlugin_setup_cacheLoad_rsp_payload_refillSlot;
  wire                MmuPlugin_setup_cacheLoad_rsp_payload_refillSlotAny;
  reg                 MmuPlugin_setup_invalidatePort_cmd_valid;
  reg                 MmuPlugin_setup_invalidatePort_rsp_valid;
  wire                FetchPlugin_stages_0_valid;
  reg                 _zz_FetchPlugin_stages_1_valid;
  reg                 FetchPlugin_stages_1_valid;
  reg                 _zz_FetchPlugin_stages_2_valid;
  reg                 FetchPlugin_stages_2_valid;
  reg                 _zz_AlignerPlugin_setup_s2m_valid;
  reg                 FetchCachePlugin_setup_redoJump_valid;
  wire       [31:0]   FetchCachePlugin_setup_redoJump_payload_pc;
  wire                FetchCachePlugin_setup_historyJump_valid;
  wire       [23:0]   FetchCachePlugin_setup_historyJump_payload_history;
  wire                FetchCachePlugin_setup_refillEvent;
  reg                 FetchCachePlugin_setup_invalidatePort_cmd_valid;
  reg                 FetchCachePlugin_setup_invalidatePort_rsp_valid;
  wire                AlignerPlugin_setup_s2m_valid;
  wire                AlignerPlugin_setup_sequenceJump_valid;
  wire       [31:0]   AlignerPlugin_setup_sequenceJump_payload_pc;
  wire                AlignerPlugin_setup_singleFetch;
  wire                FrontendPlugin_aligned_valid;
  wire                FrontendPlugin_decompressed_valid;
  wire                FrontendPlugin_decoded_valid;
  reg                 _zz_FrontendPlugin_serialized_valid;
  reg                 FrontendPlugin_serialized_valid;
  wire                _zz_FrontendPlugin_serialized_isForked;
  wire                FrontendPlugin_allocated_valid;
  reg                 _zz_FrontendPlugin_dispatch_valid;
  reg                 FrontendPlugin_dispatch_valid;
  wire                FrontendPlugin_decoded_isFireing /* verilator public */ ;
  wire                FrontendPlugin_allocated_isFireing /* verilator public */ ;
  wire                FrontendPlugin_isBusy;
  wire                FrontendPlugin_isBusyAfterDecode;
  wire                DecoderPlugin_setup_exceptionPort_valid;
  reg        [3:0]    DecoderPlugin_setup_exceptionPort_payload_cause;
  wire       [31:0]   DecoderPlugin_setup_exceptionPort_payload_epc;
  reg        [31:0]   DecoderPlugin_setup_exceptionPort_payload_tval;
  reg                 DecoderPlugin_setup_trapHalt;
  reg                 DecoderPlugin_setup_trapRaise;
  wire                DecoderPlugin_setup_trapReady;
  wire                DecoderPlugin_setup_debugEnter_0;
  wire                DecoderPlugin_setup_debugEnter_1;
  wire                BranchContextPlugin_setup_learnValid;
  wire                DecoderPredictionPlugin_setup_decodeJump_valid;
  wire       [31:0]   DecoderPredictionPlugin_setup_decodeJump_payload_pc;
  wire                DecoderPredictionPlugin_setup_historyPush_flush;
  reg        [1:0]    DecoderPredictionPlugin_setup_historyPush_mask;
  reg        [1:0]    DecoderPredictionPlugin_setup_historyPush_taken;
  reg        [23:0]   HistoryPlugin_logic_update_pushes_2_state;
  wire                BtbPlugin_setup_btbJump_valid;
  wire       [31:0]   BtbPlugin_setup_btbJump_payload_pc;
  wire                BtbPlugin_setup_historyPush_flush;
  wire       [0:0]    BtbPlugin_setup_historyPush_mask;
  wire       [0:0]    BtbPlugin_setup_historyPush_taken;
  reg        [23:0]   HistoryPlugin_logic_update_pushes_0_state;
  reg                 Lsu2Plugin_setup_postCommitBusy;
  reg        [1:0]    Lsu2Plugin_setup_fpuWriteSize;
  reg                 Lsu2Plugin_setup_regfilePorts_0_write_valid;
  reg        [5:0]    Lsu2Plugin_setup_regfilePorts_0_write_address;
  reg        [31:0]   Lsu2Plugin_setup_regfilePorts_0_write_data;
  reg        [5:0]    Lsu2Plugin_setup_regfilePorts_0_write_robId;
  reg                 Lsu2Plugin_setup_cacheLoad_cmd_valid;
  wire                Lsu2Plugin_setup_cacheLoad_cmd_ready;
  reg        [31:0]   Lsu2Plugin_setup_cacheLoad_cmd_payload_virtual;
  reg        [1:0]    Lsu2Plugin_setup_cacheLoad_cmd_payload_size;
  reg                 Lsu2Plugin_setup_cacheLoad_cmd_payload_redoOnDataHazard;
  wire                Lsu2Plugin_setup_cacheLoad_cmd_payload_unlocked;
  reg                 Lsu2Plugin_setup_cacheLoad_cmd_payload_unique;
  reg        [31:0]   Lsu2Plugin_setup_cacheLoad_translated_physical;
  reg                 Lsu2Plugin_setup_cacheLoad_translated_abord;
  wire       [2:0]    Lsu2Plugin_setup_cacheLoad_cancels;
  wire                Lsu2Plugin_setup_cacheLoad_rsp_valid;
  wire       [31:0]   Lsu2Plugin_setup_cacheLoad_rsp_payload_data;
  wire                Lsu2Plugin_setup_cacheLoad_rsp_payload_fault;
  wire                Lsu2Plugin_setup_cacheLoad_rsp_payload_redo;
  wire       [1:0]    Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlot;
  wire                Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlotAny;
  reg                 Lsu2Plugin_setup_cacheStore_cmd_valid;
  wire                Lsu2Plugin_setup_cacheStore_cmd_ready;
  reg        [31:0]   Lsu2Plugin_setup_cacheStore_cmd_payload_address;
  reg        [31:0]   Lsu2Plugin_setup_cacheStore_cmd_payload_data;
  wire       [3:0]    Lsu2Plugin_setup_cacheStore_cmd_payload_mask;
  wire                Lsu2Plugin_setup_cacheStore_cmd_payload_generation;
  reg                 Lsu2Plugin_setup_cacheStore_cmd_payload_io;
  reg                 Lsu2Plugin_setup_cacheStore_cmd_payload_flush;
  wire                Lsu2Plugin_setup_cacheStore_cmd_payload_flushFree;
  reg                 Lsu2Plugin_setup_cacheStore_cmd_payload_prefetch;
  wire                Lsu2Plugin_setup_cacheStore_rsp_valid;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_fault;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_redo;
  wire       [1:0]    Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlot;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlotAny;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_generationKo;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_flush;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_prefetch;
  wire       [31:0]   Lsu2Plugin_setup_cacheStore_rsp_payload_address;
  wire                Lsu2Plugin_setup_cacheStore_rsp_payload_io;
  reg                 Lsu2Plugin_setup_sharedCompletion_valid;
  wire       [5:0]    Lsu2Plugin_setup_sharedCompletion_payload_id;
  reg                 Lsu2Plugin_setup_sharedTrap_valid;
  reg        [5:0]    Lsu2Plugin_setup_sharedTrap_payload_robId;
  reg                 Lsu2Plugin_setup_sharedTrap_payload_trap;
  wire       [31:0]   Lsu2Plugin_setup_sharedTrap_payload_pcTarget;
  reg        [3:0]    Lsu2Plugin_setup_sharedTrap_payload_cause;
  wire       [31:0]   Lsu2Plugin_setup_sharedTrap_payload_tval;
  wire                Lsu2Plugin_setup_sharedTrap_payload_skipCommit;
  reg        [7:0]    Lsu2Plugin_setup_sharedTrap_payload_reason;
  reg                 Lsu2Plugin_setup_specialTrap_valid;
  wire       [5:0]    Lsu2Plugin_setup_specialTrap_payload_robId;
  wire       [3:0]    Lsu2Plugin_setup_specialTrap_payload_cause;
  wire       [31:0]   Lsu2Plugin_setup_specialTrap_payload_tval;
  wire                Lsu2Plugin_setup_specialTrap_payload_skipCommit;
  wire       [7:0]    Lsu2Plugin_setup_specialTrap_payload_reason;
  reg                 Lsu2Plugin_setup_specialCompletion_valid;
  wire       [5:0]    Lsu2Plugin_setup_specialCompletion_payload_id;
  reg                 Lsu2Plugin_setup_flushPort_cmd_valid;
  reg                 Lsu2Plugin_setup_flushPort_cmd_payload_withFree;
  reg                 Lsu2Plugin_setup_flushPort_rsp_valid;
  wire                DataCachePlugin_setup_writebackBusy;
  wire                DataCachePlugin_setup_refillEvent;
  wire                DataCachePlugin_setup_writebackEvent;
  wire       [1:0]    DataCachePlugin_setup_refillCompletions;
  reg                 DataCachePlugin_setup_lockPort_valid;
  reg        [31:0]   DataCachePlugin_setup_lockPort_address;
  wire                CommitPlugin_setup_jump_valid;
  wire       [31:0]   CommitPlugin_setup_jump_payload_pc;
  wire       [5:0]    CommitPlugin_setup_robLineMask_line;
  reg        [1:0]    CommitPlugin_setup_robLineMask_mask;
  wire                CommitPlugin_setup_isRobEmpty;
  reg                 PrivilegedPlugin_setup_jump_valid;
  reg        [31:0]   PrivilegedPlugin_setup_jump_payload_pc;
  reg        [1:0]    PrivilegedPlugin_setup_privilege;
  wire                PrivilegedPlugin_setup_withMachinePrivilege;
  wire                PrivilegedPlugin_setup_withSupervisorPrivilege;
  reg                 PrivilegedPlugin_setup_xretAwayFromMachine;
  reg                 PrivilegedPlugin_setup_trapEvent;
  reg                 PrivilegedPlugin_setup_redoTriggered;
  wire                PrivilegedPlugin_setup_setFpDirty;
  wire                PrivilegedPlugin_setup_isFpuEnabled;
  wire                ALU0_ExecutionUnitBase_pipeline_fetch_0_valid;
  reg                 ALU0_ExecutionUnitBase_pipeline_fetch_1_valid;
  wire                ALU0_IntAluPlugin_setup_intFormatPort_valid;
  wire       [31:0]   ALU0_IntAluPlugin_setup_intFormatPort_payload;
  wire                ALU0_ShiftPlugin_setup_intFormatPort_valid;
  wire       [31:0]   ALU0_ShiftPlugin_setup_intFormatPort_payload;
  wire                ALU0_BranchPlugin_setup_intFormatPort_valid;
  wire       [31:0]   ALU0_BranchPlugin_setup_intFormatPort_payload;
  wire                ALU0_BranchPlugin_setup_reschedule_valid;
  wire       [5:0]    ALU0_BranchPlugin_setup_reschedule_payload_robId;
  wire                ALU0_BranchPlugin_setup_reschedule_payload_trap;
  wire       [31:0]   ALU0_BranchPlugin_setup_reschedule_payload_pcTarget;
  wire       [3:0]    ALU0_BranchPlugin_setup_reschedule_payload_cause;
  wire       [31:0]   ALU0_BranchPlugin_setup_reschedule_payload_tval;
  wire                ALU0_BranchPlugin_setup_reschedule_payload_skipCommit;
  wire       [7:0]    ALU0_BranchPlugin_setup_reschedule_payload_reason;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_0_valid;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_1_valid;
  wire                EU0_MulPlugin_setup_intFormatPort_valid;
  wire       [31:0]   EU0_MulPlugin_setup_intFormatPort_payload;
  wire                EU0_DivPlugin_setup_intFormatPort_valid;
  wire       [31:0]   EU0_DivPlugin_setup_intFormatPort_payload;
  wire                AguPlugin_setup_port_valid /* verilator public */ ;
  wire       [5:0]    AguPlugin_setup_port_payload_robId /* verilator public */ ;
  wire       [0:0]    AguPlugin_setup_port_payload_robIdMsb;
  wire       [4:0]    AguPlugin_setup_port_payload_aguId /* verilator public */ ;
  wire                AguPlugin_setup_port_payload_load /* verilator public */ ;
  wire       [31:0]   AguPlugin_setup_port_payload_address;
  wire       [1:0]    AguPlugin_setup_port_payload_size;
  wire                AguPlugin_setup_port_payload_unsigned;
  wire       [5:0]    AguPlugin_setup_port_payload_physicalRd;
  wire                AguPlugin_setup_port_payload_writeRd;
  wire       [31:0]   AguPlugin_setup_port_payload_pc;
  wire                AguPlugin_setup_port_payload_lr;
  wire                AguPlugin_setup_port_payload_earlySample;
  wire       [31:0]   AguPlugin_setup_port_payload_earlyPc;
  wire       [31:0]   AguPlugin_setup_port_payload_data /* verilator public */ ;
  wire                AguPlugin_setup_port_payload_amo;
  wire                AguPlugin_setup_port_payload_sc;
  wire                AguPlugin_setup_port_payload_swap;
  wire       [2:0]    AguPlugin_setup_port_payload_op;
  wire                EnvCallPlugin_setup_reschedule_valid;
  wire       [5:0]    EnvCallPlugin_setup_reschedule_payload_robId;
  reg        [3:0]    EnvCallPlugin_setup_reschedule_payload_cause;
  reg        [31:0]   EnvCallPlugin_setup_reschedule_payload_tval;
  reg                 EnvCallPlugin_setup_reschedule_payload_skipCommit;
  reg        [7:0]    EnvCallPlugin_setup_reschedule_payload_reason;
  wire                EU0_CsrAccessPlugin_setup_intFormatPort_valid;
  wire       [31:0]   EU0_CsrAccessPlugin_setup_intFormatPort_payload;
  reg                 EU0_CsrAccessPlugin_setup_onDecodeTrap;
  reg                 EU0_CsrAccessPlugin_setup_onDecodeFlushPipeline;
  wire                EU0_CsrAccessPlugin_setup_onDecodeRead;
  wire                EU0_CsrAccessPlugin_setup_onDecodeWrite;
  wire       [11:0]   EU0_CsrAccessPlugin_setup_onDecodeAddress;
  reg                 EU0_CsrAccessPlugin_setup_onReadHalt;
  reg                 EU0_CsrAccessPlugin_setup_onWriteHalt;
  reg        [31:0]   EU0_CsrAccessPlugin_setup_onReadToWriteBits;
  wire       [31:0]   EU0_CsrAccessPlugin_setup_onWriteBits;
  wire       [11:0]   EU0_CsrAccessPlugin_setup_onWriteAddress;
  wire                EU0_CsrAccessPlugin_setup_onWriteFlushPipeline;
  wire       [11:0]   EU0_CsrAccessPlugin_setup_onReadAddress;
  wire                EU0_CsrAccessPlugin_setup_onReadMovingOff;
  wire                EU0_CsrAccessPlugin_setup_onWriteMovingOff;
  wire                EU0_CsrAccessPlugin_setup_trap_valid;
  wire       [5:0]    EU0_CsrAccessPlugin_setup_trap_payload_robId;
  reg        [3:0]    EU0_CsrAccessPlugin_setup_trap_payload_cause;
  wire       [31:0]   EU0_CsrAccessPlugin_setup_trap_payload_tval;
  wire                EU0_CsrAccessPlugin_setup_trap_payload_skipCommit;
  wire       [7:0]    EU0_CsrAccessPlugin_setup_trap_payload_reason;
  wire                ALU1_ExecutionUnitBase_pipeline_fetch_0_valid;
  reg                 ALU1_ExecutionUnitBase_pipeline_fetch_1_valid;
  wire                ALU1_IntAluPlugin_setup_intFormatPort_valid;
  wire       [31:0]   ALU1_IntAluPlugin_setup_intFormatPort_payload;
  wire                ALU1_ShiftPlugin_setup_intFormatPort_valid;
  wire       [31:0]   ALU1_ShiftPlugin_setup_intFormatPort_payload;
  wire                ALU1_BranchPlugin_setup_intFormatPort_valid;
  wire       [31:0]   ALU1_BranchPlugin_setup_intFormatPort_payload;
  wire                ALU1_BranchPlugin_setup_reschedule_valid;
  wire       [5:0]    ALU1_BranchPlugin_setup_reschedule_payload_robId;
  wire                ALU1_BranchPlugin_setup_reschedule_payload_trap;
  wire       [31:0]   ALU1_BranchPlugin_setup_reschedule_payload_pcTarget;
  wire       [3:0]    ALU1_BranchPlugin_setup_reschedule_payload_cause;
  wire       [31:0]   ALU1_BranchPlugin_setup_reschedule_payload_tval;
  wire                ALU1_BranchPlugin_setup_reschedule_payload_skipCommit;
  wire       [7:0]    ALU1_BranchPlugin_setup_reschedule_payload_reason;
  wire                FetchPlugin_stages_1_isFireing;
  reg                 _zz_FetchPlugin_stages_1_isFirstCycle;
  wire                when_Stage_l170;
  wire                FetchPlugin_stages_1_isFirstCycle /* verilator public */ ;
  wire       [5:0]    _zz_PcPlugin_logic_jump_oh;
  wire                _zz_PcPlugin_logic_jump_oh_1;
  wire                _zz_PcPlugin_logic_jump_oh_2;
  wire                _zz_PcPlugin_logic_jump_oh_3;
  wire                _zz_PcPlugin_logic_jump_oh_4;
  wire                _zz_PcPlugin_logic_jump_oh_5;
  reg        [5:0]    _zz_PcPlugin_logic_jump_oh_6;
  wire       [5:0]    PcPlugin_logic_jump_oh;
  (* keep , syn_keep *) wire       [31:0]   PcPlugin_logic_jump_target /* synthesis syn_keep = 1 */ ;
  wire                _zz_PcPlugin_logic_jump_target_1;
  wire                when_PcPlugin_l55;
  wire                PcPlugin_logic_jump_pcLoad_valid;
  wire       [31:0]   PcPlugin_logic_jump_pcLoad_payload_pc;
  wire                FetchCachePlugin_logic_translationPort_wake;
  wire                FetchCachePlugin_logic_banks_0_write_valid;
  wire       [8:0]    FetchCachePlugin_logic_banks_0_write_payload_address;
  wire       [63:0]   FetchCachePlugin_logic_banks_0_write_payload_data;
  wire                FetchCachePlugin_logic_banks_0_read_cmd_valid;
  wire       [8:0]    FetchCachePlugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchCachePlugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                FetchCachePlugin_logic_banks_1_write_valid;
  wire       [8:0]    FetchCachePlugin_logic_banks_1_write_payload_address;
  wire       [63:0]   FetchCachePlugin_logic_banks_1_write_payload_data;
  wire                FetchCachePlugin_logic_banks_1_read_cmd_valid;
  wire       [8:0]    FetchCachePlugin_logic_banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchCachePlugin_logic_banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                FetchCachePlugin_logic_banks_2_write_valid;
  wire       [8:0]    FetchCachePlugin_logic_banks_2_write_payload_address;
  wire       [63:0]   FetchCachePlugin_logic_banks_2_write_payload_data;
  wire                FetchCachePlugin_logic_banks_2_read_cmd_valid;
  wire       [8:0]    FetchCachePlugin_logic_banks_2_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchCachePlugin_logic_banks_2_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                FetchCachePlugin_logic_banks_3_write_valid;
  wire       [8:0]    FetchCachePlugin_logic_banks_3_write_payload_address;
  wire       [63:0]   FetchCachePlugin_logic_banks_3_write_payload_data;
  wire                FetchCachePlugin_logic_banks_3_read_cmd_valid;
  wire       [8:0]    FetchCachePlugin_logic_banks_3_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchCachePlugin_logic_banks_3_read_rsp /* synthesis syn_keep = 1 */ ;
  reg        [3:0]    FetchCachePlugin_logic_waysWrite_mask;
  reg        [5:0]    FetchCachePlugin_logic_waysWrite_address;
  reg                 FetchCachePlugin_logic_waysWrite_tag_loaded;
  reg                 FetchCachePlugin_logic_waysWrite_tag_error;
  reg        [19:0]   FetchCachePlugin_logic_waysWrite_tag_address;
  wire                FetchCachePlugin_logic_ways_0_read_cmd_valid;
  wire       [5:0]    FetchCachePlugin_logic_ways_0_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_0_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_0_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchCachePlugin_logic_ways_0_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded;
  wire                FetchCachePlugin_logic_ways_1_read_cmd_valid;
  wire       [5:0]    FetchCachePlugin_logic_ways_1_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_1_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_1_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchCachePlugin_logic_ways_1_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_1_read_rsp_loaded;
  wire                FetchCachePlugin_logic_ways_2_read_cmd_valid;
  wire       [5:0]    FetchCachePlugin_logic_ways_2_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_2_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_2_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchCachePlugin_logic_ways_2_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_2_read_rsp_loaded;
  wire                FetchCachePlugin_logic_ways_3_read_cmd_valid;
  wire       [5:0]    FetchCachePlugin_logic_ways_3_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_3_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchCachePlugin_logic_ways_3_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchCachePlugin_logic_ways_3_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchCachePlugin_logic_ways_3_read_rsp_loaded;
  reg                 FetchCachePlugin_logic_plru_write_valid;
  reg        [5:0]    FetchCachePlugin_logic_plru_write_payload_address;
  reg        [0:0]    FetchCachePlugin_logic_plru_write_payload_data_0;
  reg        [1:0]    FetchCachePlugin_logic_plru_write_payload_data_1;
  reg                 FetchCachePlugin_logic_invalidate_requested;
  reg                 FetchCachePlugin_logic_invalidate_canStart;
  reg        [6:0]    FetchCachePlugin_logic_invalidate_counter;
  wire                FetchCachePlugin_logic_invalidate_done;
  reg                 FetchCachePlugin_logic_invalidate_firstEver;
  wire                when_FetchCachePlugin_l379;
  wire                when_FetchCachePlugin_l383;
  wire                FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l389;
  wire                when_FetchCachePlugin_l391;
  wire                when_FetchCachePlugin_l396;
  reg                 FetchCachePlugin_logic_invalidate_done_regNext;
  wire                when_FetchCachePlugin_l400;
  reg                 FetchCachePlugin_logic_refill_start_valid;
  wire       [31:0]   FetchCachePlugin_logic_refill_start_address;
  wire       [1:0]    FetchCachePlugin_logic_refill_start_wayToAllocate;
  wire                FetchCachePlugin_logic_refill_start_isIo;
  reg                 FetchCachePlugin_logic_refill_fire;
  reg                 FetchCachePlugin_logic_refill_valid;
  (* keep , syn_keep *) reg        [31:0]   FetchCachePlugin_logic_refill_address /* synthesis syn_keep = 1 */ ;
  reg                 FetchCachePlugin_logic_refill_isIo;
  reg                 FetchCachePlugin_logic_refill_hadError;
  reg        [1:0]    FetchCachePlugin_logic_refill_wayToAllocate;
  reg        [31:0]   FetchCachePlugin_logic_refill_pushCounter;
  wire                when_FetchCachePlugin_l422;
  reg                 FetchCachePlugin_logic_refill_cmdSent;
  wire                FetchCachePlugin_mem_cmd_fire;
  wire                when_Utils_l560;
  reg                 FetchCachePlugin_logic_refill_randomWay_willIncrement;
  wire                FetchCachePlugin_logic_refill_randomWay_willClear;
  reg        [1:0]    FetchCachePlugin_logic_refill_randomWay_valueNext;
  reg        [1:0]    FetchCachePlugin_logic_refill_randomWay_value;
  wire                FetchCachePlugin_logic_refill_randomWay_willOverflowIfInc;
  wire                FetchCachePlugin_logic_refill_randomWay_willOverflow;
  (* keep , syn_keep *) reg        [2:0]    FetchCachePlugin_logic_refill_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                when_FetchCachePlugin_l470;
  wire                FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l476;
  reg                 FetchCachePlugin_logic_refill_fire_regNext;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_0;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_1;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_2;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_3;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_4;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_5;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_translatedHits;
  wire                FetchCachePlugin_logic_read_onWays_0_hits_bypassHits;
  wire                FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_0;
  wire                FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_1;
  wire                FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_2;
  wire                FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_3;
  wire                FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_4;
  wire                FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_5;
  wire                FetchCachePlugin_logic_read_onWays_1_hits_translatedHits;
  wire                FetchCachePlugin_logic_read_onWays_1_hits_bypassHits;
  wire                FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_0;
  wire                FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_1;
  wire                FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_2;
  wire                FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_3;
  wire                FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_4;
  wire                FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_5;
  wire                FetchCachePlugin_logic_read_onWays_2_hits_translatedHits;
  wire                FetchCachePlugin_logic_read_onWays_2_hits_bypassHits;
  wire                FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_0;
  wire                FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_1;
  wire                FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_2;
  wire                FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_3;
  wire                FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_4;
  wire                FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_5;
  wire                FetchCachePlugin_logic_read_onWays_3_hits_translatedHits;
  wire                FetchCachePlugin_logic_read_onWays_3_hits_bypassHits;
  wire       [5:0]    _zz_FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0;
  wire       [2:0]    _zz_FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0_1;
  wire       [0:0]    FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_context_state_0;
  wire       [1:0]    FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_context_state_1;
  wire       [1:0]    FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_evict_id;
  wire       [1:0]    FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_state_0;
  reg        [1:0]    FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_state_1;
  wire                FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_sel_0;
  wire                FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_sel_1;
  wire                FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_logic_0_state;
  wire       [0:0]    FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_logic_1_stateSel;
  wire                FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_logic_1_state;
  wire       [0:0]    FetchCachePlugin_logic_read_ctrl_plruLogic_core_update_logic_1_sel;
  wire                _zz_FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id;
  wire                _zz_FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id_1;
  reg                 FetchCachePlugin_logic_read_ctrl_redoIt;
  wire                FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552;
  wire                FetchPlugin_stages_2_isFireing;
  wire                when_FetchCachePlugin_l562;
  wire                FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l583;
  wire                when_FetchCachePlugin_l593;
  wire       [2:0]    _zz_FetchCachePlugin_logic_plru_write_payload_data_0;
  wire                AlignerPlugin_logic_ignoreInput;
  wire                AlignerPlugin_logic_isInputValid;
  wire                when_AlignerPlugin_l98;
  reg        [63:0]   AlignerPlugin_logic_buffer_data;
  reg        [1:0]    AlignerPlugin_logic_buffer_mask;
  reg        [31:0]   AlignerPlugin_logic_buffer_pc;
  reg                 AlignerPlugin_logic_buffer_fault;
  reg                 AlignerPlugin_logic_buffer_fault_page;
  reg                 AlignerPlugin_logic_buffer_branchValid;
  reg        [0:0]    AlignerPlugin_logic_buffer_branchSlice;
  reg        [31:0]   AlignerPlugin_logic_buffer_branchPcNext;
  reg        [23:0]   AlignerPlugin_logic_buffer_wordContexts_0;
  reg                 AlignerPlugin_logic_buffer_wordContexts_1;
  reg        [0:0]    AlignerPlugin_logic_buffer_wordContexts_2;
  reg                 AlignerPlugin_logic_buffer_wordContexts_3;
  reg        [1:0]    AlignerPlugin_logic_buffer_wordContexts_4_0;
  reg        [1:0]    AlignerPlugin_logic_buffer_wordContexts_4_1;
  reg        [11:0]   AlignerPlugin_logic_buffer_firstWordContexts_0;
  wire       [127:0]  _zz_AlignerPlugin_logic_slices_data_0;
  wire       [31:0]   AlignerPlugin_logic_slices_data_0;
  wire       [31:0]   AlignerPlugin_logic_slices_data_1;
  wire       [31:0]   AlignerPlugin_logic_slices_data_2;
  wire       [31:0]   AlignerPlugin_logic_slices_data_3;
  wire       [3:0]    AlignerPlugin_logic_slices_carry;
  wire       [3:0]    AlignerPlugin_logic_slices_remains;
  wire       [3:0]    AlignerPlugin_logic_slices_used;
  wire       [3:0]    AlignerPlugin_logic_decoders_0_usage;
  wire                AlignerPlugin_logic_decoders_0_notEnoughData;
  wire                AlignerPlugin_logic_decoders_0_pastPrediction;
  wire                AlignerPlugin_logic_decoders_0_usable;
  wire       [3:0]    AlignerPlugin_logic_decoders_1_usage;
  wire                AlignerPlugin_logic_decoders_1_notEnoughData;
  wire                AlignerPlugin_logic_decoders_1_pastPrediction;
  wire                AlignerPlugin_logic_decoders_1_usable;
  wire       [3:0]    AlignerPlugin_logic_decoders_2_usage;
  wire                AlignerPlugin_logic_decoders_2_notEnoughData;
  wire                AlignerPlugin_logic_decoders_2_pastPrediction;
  wire                AlignerPlugin_logic_decoders_2_usable;
  wire       [3:0]    AlignerPlugin_logic_decoders_3_usage;
  wire                AlignerPlugin_logic_decoders_3_notEnoughData;
  wire                AlignerPlugin_logic_decoders_3_pastPrediction;
  wire                AlignerPlugin_logic_decoders_3_usable;
  wire                _zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1;
  wire       [3:0]    _zz_AlignerPlugin_logic_extractors_0_maskOh;
  wire                _zz_AlignerPlugin_logic_extractors_0_maskOh_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_maskOh_2;
  wire                _zz_AlignerPlugin_logic_extractors_0_maskOh_3;
  reg        [3:0]    _zz_AlignerPlugin_logic_extractors_0_maskOh_4;
  wire       [3:0]    AlignerPlugin_logic_extractors_0_maskOh;
  wire                _zz_AlignerPlugin_logic_extractors_0_usage;
  wire                _zz_AlignerPlugin_logic_extractors_0_usage_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_usage_2;
  wire                _zz_AlignerPlugin_logic_extractors_0_usage_3;
  wire       [3:0]    AlignerPlugin_logic_extractors_0_usage;
  wire                AlignerPlugin_logic_extractors_0_usable;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_slice0;
  wire                AlignerPlugin_logic_extractors_0_valid;
  wire       [0:0]    AlignerPlugin_logic_extractors_0_sliceLast;
  wire                AlignerPlugin_logic_extractors_0_bufferPredictionLast;
  wire                AlignerPlugin_logic_extractors_0_inputPredictionLast;
  wire                AlignerPlugin_logic_extractors_0_lastWord;
  wire       [3:0]    _zz_AlignerPlugin_logic_extractors_0_sliceOffset;
  wire                _zz_AlignerPlugin_logic_extractors_0_sliceOffset_1;
  wire                _zz_AlignerPlugin_logic_extractors_0_sliceOffset_2;
  wire                _zz_AlignerPlugin_logic_extractors_0_sliceOffset_3;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_sliceOffset;
  wire                AlignerPlugin_logic_extractors_0_firstWord;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_pcWord;
  wire                when_AlignerPlugin_l230;
  wire                when_AlignerPlugin_l235;
  wire       [2:0]    _zz_AlignerPlugin_logic_extractors_1_maskOh;
  wire                _zz_AlignerPlugin_logic_extractors_1_maskOh_1;
  wire                _zz_AlignerPlugin_logic_extractors_1_maskOh_2;
  reg        [2:0]    _zz_AlignerPlugin_logic_extractors_1_maskOh_3;
  wire       [2:0]    AlignerPlugin_logic_extractors_1_maskOh;
  wire                _zz_AlignerPlugin_logic_extractors_1_usage;
  wire                _zz_AlignerPlugin_logic_extractors_1_usage_1;
  wire                _zz_AlignerPlugin_logic_extractors_1_usage_2;
  wire       [3:0]    AlignerPlugin_logic_extractors_1_usage;
  wire                AlignerPlugin_logic_extractors_1_usable;
  wire       [31:0]   AlignerPlugin_logic_extractors_1_slice0;
  reg                 AlignerPlugin_logic_extractors_1_valid;
  wire       [0:0]    AlignerPlugin_logic_extractors_1_sliceLast;
  wire                AlignerPlugin_logic_extractors_1_bufferPredictionLast;
  wire                AlignerPlugin_logic_extractors_1_inputPredictionLast;
  wire                AlignerPlugin_logic_extractors_1_lastWord;
  wire       [3:0]    _zz_AlignerPlugin_logic_extractors_1_sliceOffset;
  wire                _zz_AlignerPlugin_logic_extractors_1_sliceOffset_1;
  wire                _zz_AlignerPlugin_logic_extractors_1_sliceOffset_2;
  wire                _zz_AlignerPlugin_logic_extractors_1_sliceOffset_3;
  wire       [1:0]    AlignerPlugin_logic_extractors_1_sliceOffset;
  wire                AlignerPlugin_logic_extractors_1_firstWord;
  wire       [31:0]   AlignerPlugin_logic_extractors_1_pcWord;
  wire                when_AlignerPlugin_l230_1;
  wire                when_AlignerPlugin_l235_1;
  wire                FrontendPlugin_aligned_isFireing;
  wire                AlignerPlugin_logic_fireOutput;
  wire                AlignerPlugin_logic_fireInput;
  wire       [1:0]    AlignerPlugin_logic_postMask;
  reg                 AlignerPlugin_logic_correctionSent;
  wire                when_AlignerPlugin_l264;
  wire                _zz_FetchPlugin_stages_1_isFlushingRoot;
  wire                AlignerPlugin_setup_s2m_haltRequest_AlignerPlugin_l270;
  wire                integer_RfAllocationPlugin_logic_pop_blocked;
  wire                FrontendPlugin_allocated_haltRequest_RfAllocationPlugin_l55;
  wire                when_RfAllocationPlugin_l63;
  wire                when_RfAllocationPlugin_l63_1;
  reg        [1:0]    DispatchPlugin_logic_sparseRob_todo;
  wire       [1:0]    DispatchPlugin_logic_sparseRob_mask;
  wire       [1:0]    DispatchPlugin_logic_sparseRob_remains;
  wire       [1:0]    DispatchPlugin_logic_sparseRob_sparse;
  wire                DispatchPlugin_logic_sparseRob_sparseHit;
  wire       [1:0]    DispatchPlugin_logic_sparseRob_sparse_ohFirst_input;
  wire       [1:0]    DispatchPlugin_logic_sparseRob_sparse_ohFirst_masked;
  wire       [1:0]    DispatchPlugin_logic_sparseRob_sparseFirst;
  reg        [1:0]    DispatchPlugin_logic_sparseRob_filter;
  wire                when_DispatchPlugin_l79;
  wire                when_DispatchPlugin_l79_1;
  wire       [1:0]    DispatchPlugin_logic_sparseRob_masked;
  wire                DispatchPlugin_logic_sparseRob_forkLast;
  wire                FrontendPlugin_serialized_forkRequest_DispatchPlugin_l90;
  wire                when_DispatchPlugin_l94;
  reg        [4:0]    BranchContextPlugin_logic_ptr_alloc;
  reg        [4:0]    BranchContextPlugin_logic_ptr_commited;
  reg        [4:0]    BranchContextPlugin_logic_ptr_free;
  wire       [4:0]    BranchContextPlugin_logic_ptr_occupancy;
  wire       [4:0]    BranchContextPlugin_logic_alloc_allocNext;
  reg                 BranchContextPlugin_logic_alloc_full;
  wire                when_BranchContextPlugin_l93;
  wire                when_BranchContextPlugin_l93_1;
  wire                when_BranchContextPlugin_l106;
  wire                FrontendPlugin_allocated_haltRequest_BranchContextPlugin_l107;
  reg        [23:0]   HistoryPlugin_logic_onCommit_value /* verilator public */ ;
  wire       [23:0]   HistoryPlugin_logic_onCommit_whitebox_0 /* verilator public */ ;
  wire       [23:0]   HistoryPlugin_logic_onCommit_whitebox_1 /* verilator public */ ;
  reg        [3:0]    DecoderPredictionPlugin_logic_ras_ptr_push;
  reg        [3:0]    DecoderPredictionPlugin_logic_ras_ptr_pop;
  reg                 DecoderPredictionPlugin_logic_ras_ptr_pushIt;
  reg                 DecoderPredictionPlugin_logic_ras_ptr_popIt;
  wire       [31:0]   DecoderPredictionPlugin_logic_ras_read;
  wire                DecoderPredictionPlugin_logic_ras_write_valid;
  wire       [3:0]    DecoderPredictionPlugin_logic_ras_write_payload_address;
  reg        [31:0]   DecoderPredictionPlugin_logic_ras_write_payload_data;
  wire       [31:0]   BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice;
  wire       [31:0]   BranchContextPlugin_learn_BRANCH_FINAL_pcTarget;
  wire                BranchContextPlugin_learn_BRANCH_FINAL_taken;
  wire       [15:0]   BtbPlugin_logic_onLearn_hash;
  wire                BtbPlugin_logic_onLearn_port_valid;
  wire       [8:0]    BtbPlugin_logic_onLearn_port_payload_address;
  wire       [15:0]   BtbPlugin_logic_onLearn_port_payload_data_hash;
  wire       [0:0]    BtbPlugin_logic_onLearn_port_payload_data_slice;
  wire       [31:0]   BtbPlugin_logic_onLearn_port_payload_data_pcTarget;
  wire                BtbPlugin_logic_onLearn_port_payload_data_isBranch;
  wire                BranchContextPlugin_free_learn_Prediction_IS_BRANCH;
  wire       [8:0]    BtbPlugin_logic_readCmd_entryAddress;
  wire       [49:0]   _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash;
  wire                BtbPlugin_logic_hitCalc_postPcPrediction;
  wire                BtbPlugin_logic_applyIt_prediction;
  wire                BtbPlugin_logic_applyIt_needIt;
  reg                 BtbPlugin_logic_applyIt_correctionSent;
  wire                when_BtbPlugin_l109;
  wire                BtbPlugin_logic_applyIt_doIt;
  wire                GSharePlugin_logic_mem_write_valid;
  wire       [12:0]   GSharePlugin_logic_mem_write_payload_address;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_0;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_1;
  wire       [12:0]   _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH;
  wire       [3:0]    _zz_FetchPlugin_stages_1_GSHARE_COUNTER_0;
  wire                when_GSharePlugin_l98;
  wire       [23:0]   BranchContextPlugin_free_learn_BRANCH_HISTORY;
  wire       [12:0]   _zz_GSharePlugin_logic_onLearn_hash;
  wire       [12:0]   GSharePlugin_logic_onLearn_hash;
  wire       [1:0]    BranchContextPlugin_free_learn_GSHARE_COUNTER_0;
  wire       [1:0]    BranchContextPlugin_free_learn_GSHARE_COUNTER_1;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_0;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_1;
  wire       [1:0]    GSharePlugin_logic_onLearn_incrValue;
  reg                 GSharePlugin_logic_onLearn_overflow;
  wire                when_GSharePlugin_l123;
  wire                when_GSharePlugin_l123_1;
  reg                 toplevel_DataCachePlugin_logic_cache_io_refillEvent_regNext;
  reg                 toplevel_DataCachePlugin_logic_cache_io_writebackEvent_regNext;
  wire       [1:0]    DataCachePlugin_logic_load_hits;
  wire                DataCachePlugin_logic_load_hit;
  wire       [1:0]    _zz_DataCachePlugin_logic_load_hits_bools_0;
  wire                DataCachePlugin_logic_load_hits_bools_0;
  wire                DataCachePlugin_logic_load_hits_bools_1;
  reg        [1:0]    _zz_DataCachePlugin_logic_load_oh;
  wire       [1:0]    DataCachePlugin_logic_load_oh;
  wire       [1:0]    DataCachePlugin_logic_load_ohHistory_0;
  wire       [1:0]    DataCachePlugin_logic_load_ohHistory_1;
  wire       [1:0]    DataCachePlugin_logic_load_ohHistory_2;
  wire       [1:0]    _zz_DataCachePlugin_logic_load_ohHistory_0;
  reg        [1:0]    _zz_DataCachePlugin_logic_load_ohHistory_1;
  reg        [1:0]    _zz_DataCachePlugin_logic_load_ohHistory_2;
  wire                _zz_MmuPlugin_setup_cacheLoad_cmd_ready;
  wire                _zz_io_load_translated_physical;
  reg        [6:0]    CommitPlugin_logic_ptr_alloc;
  reg        [6:0]    CommitPlugin_logic_ptr_commit;
  reg        [6:0]    CommitPlugin_logic_ptr_free;
  wire       [5:0]    CommitPlugin_logic_ptr_commitRow;
  reg        [6:0]    CommitPlugin_logic_ptr_commitNext;
  wire       [6:0]    CommitPlugin_logic_ptr_allocNext;
  wire                CommitPlugin_logic_ptr_full;
  reg                 CommitPlugin_logic_ptr_empty;
  wire                CommitPlugin_logic_ptr_canFree;
  reg        [1:0]    CommitPlugin_logic_ptr_robLineMaskRsp;
  wire                FrontendPlugin_allocated_haltRequest_CommitPlugin_l95;
  reg                 CommitPlugin_logic_reschedule_fresh;
  reg                 CommitPlugin_logic_reschedule_valid;
  reg                 CommitPlugin_logic_reschedule_trap;
  reg                 CommitPlugin_logic_reschedule_skipCommit;
  reg        [5:0]    CommitPlugin_logic_reschedule_robId;
  reg        [31:0]   CommitPlugin_logic_reschedule_pcTarget;
  reg        [3:0]    CommitPlugin_logic_reschedule_cause;
  reg        [31:0]   CommitPlugin_logic_reschedule_tval;
  reg        [7:0]    CommitPlugin_logic_reschedule_reason;
  wire       [4:0]    CommitPlugin_logic_reschedule_commit_row;
  wire       [0:0]    CommitPlugin_logic_reschedule_commit_col;
  wire                CommitPlugin_logic_reschedule_commit_rowHit;
  wire       [5:0]    CommitPlugin_logic_reschedule_age;
  wire       [5:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_0_age;
  wire       [5:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_1_age;
  wire       [5:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_2_age;
  wire       [5:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_3_age;
  wire       [5:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_4_age;
  wire       [5:0]    CommitPlugin_logic_reschedule_portsLogic_perPort_5_age;
  reg        [5:0]    CommitPlugin_logic_reschedule_portsLogic_hits;
  wire                when_CommitPlugin_l131;
  wire                _zz_CommitPlugin_logic_reschedule_trap;
  wire                _zz_CommitPlugin_logic_reschedule_trap_1;
  wire                _zz_CommitPlugin_logic_reschedule_trap_2;
  wire                _zz_CommitPlugin_logic_reschedule_trap_3;
  wire                _zz_CommitPlugin_logic_reschedule_trap_4;
  wire                _zz_CommitPlugin_logic_reschedule_trap_5;
  wire                CommitPlugin_logic_reschedule_reschedulePort_valid;
  wire       [5:0]    CommitPlugin_logic_reschedule_reschedulePort_payload_robId;
  wire                CommitPlugin_logic_reschedule_reschedulePort_payload_trap;
  wire       [3:0]    CommitPlugin_logic_reschedule_reschedulePort_payload_cause;
  wire       [31:0]   CommitPlugin_logic_reschedule_reschedulePort_payload_tval;
  wire       [7:0]    CommitPlugin_logic_reschedule_reschedulePort_payload_reason;
  wire                CommitPlugin_logic_reschedule_reschedulePort_payload_skipCommit;
  reg                 CommitPlugin_logic_commit_rescheduleHit;
  wire       [1:0]    CommitPlugin_logic_commit_active;
  reg        [1:0]    CommitPlugin_logic_commit_mask;
  reg        [1:0]    CommitPlugin_logic_commit_maskComb;
  wire                CommitPlugin_logic_commit_lineCommited;
  wire       [5:0]    CommitPlugin_logic_commit_event_robId;
  reg        [1:0]    CommitPlugin_logic_commit_event_mask;
  reg                 CommitPlugin_logic_commit_lineEvent_valid;
  wire       [5:0]    CommitPlugin_logic_commit_lineEvent_payload_robId;
  wire       [1:0]    CommitPlugin_logic_commit_lineEvent_payload_mask;
  wire                CommitPlugin_logic_commit_reschedulePort_valid;
  wire       [5:0]    CommitPlugin_logic_commit_reschedulePort_payload_robId;
  wire       [5:0]    CommitPlugin_logic_commit_reschedulePort_payload_robIdNext;
  wire                CommitPlugin_logic_commit_reschedulePort_payload_trap;
  wire       [3:0]    CommitPlugin_logic_commit_reschedulePort_payload_cause;
  wire       [31:0]   CommitPlugin_logic_commit_reschedulePort_payload_tval;
  wire       [7:0]    CommitPlugin_logic_commit_reschedulePort_payload_reason;
  wire                CommitPlugin_logic_commit_reschedulePort_payload_skipCommit;
  wire       [5:0]    CommitPlugin_logic_commit_head;
  reg        [5:0]    CommitPlugin_logic_commit_headNext;
  wire       [1:0]    _zz_CommitPlugin_logic_commit_head;
  wire                _zz_CommitPlugin_logic_commit_head_1;
  wire                CommitPlugin_logic_commit_continue;
  wire                when_CommitPlugin_l194;
  wire                CommitPlugin_commit_slot_0_enable;
  wire                CommitPlugin_commit_slot_0_readyForCommit;
  wire                CommitPlugin_commit_slot_0_rescheduleHitSlot;
  wire                when_CommitPlugin_l203;
  wire                when_CommitPlugin_l207;
  wire                when_CommitPlugin_l211;
  wire                CommitPlugin_commit_slot_1_enable;
  wire                CommitPlugin_commit_slot_1_readyForCommit;
  wire                CommitPlugin_commit_slot_1_rescheduleHitSlot;
  wire                when_CommitPlugin_l203_1;
  wire                when_CommitPlugin_l207_1;
  wire                when_CommitPlugin_l211_1;
  wire                when_CommitPlugin_l217;
  wire                CommitPlugin_logic_free_lineEventStream_valid;
  wire                CommitPlugin_logic_free_lineEventStream_ready;
  wire       [5:0]    CommitPlugin_logic_free_lineEventStream_payload_robId;
  wire       [1:0]    CommitPlugin_logic_free_lineEventStream_payload_mask;
  wire                CommitPlugin_logic_free_robHit;
  wire                CommitPlugin_logic_free_hit;
  wire                CommitPlugin_logic_free_port_valid;
  wire       [5:0]    CommitPlugin_logic_free_port_payload_robId;
  wire       [1:0]    CommitPlugin_logic_free_port_payload_commited;
  wire                robToPc_valid /* verilator public */ ;
  wire       [5:0]    robToPc_robId /* verilator public */ ;
  wire       [31:0]   robToPc_pc_0 /* verilator public */ ;
  wire       [31:0]   robToPc_pc_1 /* verilator public */ ;
  wire       [5:0]    commit_robId /* verilator public */ ;
  wire       [1:0]    commit_mask /* verilator public */ ;
  wire                reschedule_valid /* verilator public */ ;
  wire       [5:0]    reschedule_payload_robId /* verilator public */ ;
  wire       [5:0]    reschedule_payload_robIdNext /* verilator public */ ;
  wire                reschedule_payload_trap /* verilator public */ ;
  wire       [3:0]    reschedule_payload_cause /* verilator public */ ;
  wire       [31:0]   reschedule_payload_tval /* verilator public */ ;
  wire       [7:0]    reschedule_payload_reason /* verilator public */ ;
  wire                reschedule_payload_skipCommit /* verilator public */ ;
  wire       [7:0]    rescheduleReason /* verilator public */ ;
  wire       [31:0]   commit_pc_0 /* verilator public */ ;
  wire       [31:0]   commit_pc_1 /* verilator public */ ;
  wire                _zz_CommitDebugFilterPlugin_logic_commits;
  wire                _zz_CommitDebugFilterPlugin_logic_commits_1;
  wire       [17:0]   CommitDebugFilterPlugin_logic_commits;
  reg        [31:0]   CommitDebugFilterPlugin_logic_filters_0_value;
  reg        [31:0]   CommitDebugFilterPlugin_logic_filters_1_value;
  reg        [31:0]   CommitDebugFilterPlugin_logic_filters_2_value;
  wire       [1:0]    PrivilegedPlugin_logic_defaultTrap_csrPrivilege;
  wire                PrivilegedPlugin_logic_defaultTrap_csrReadOnly;
  wire                when_PrivilegedPlugin_l165;
  reg                 PrivilegedPlugin_logic_machine_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_machine_cause_code;
  reg                 PrivilegedPlugin_logic_machine_mstatus_mie;
  reg                 PrivilegedPlugin_logic_machine_mstatus_mpie;
  reg        [1:0]    PrivilegedPlugin_logic_machine_mstatus_mpp;
  reg        [1:0]    PrivilegedPlugin_logic_machine_mstatus_fs;
  reg                 PrivilegedPlugin_logic_machine_mstatus_sd;
  wire                when_PrivilegedPlugin_l393;
  reg                 PrivilegedPlugin_logic_machine_mip_meip;
  reg                 PrivilegedPlugin_logic_machine_mip_mtip;
  reg                 PrivilegedPlugin_logic_machine_mip_msip;
  reg                 PrivilegedPlugin_logic_machine_mie_meie;
  reg                 PrivilegedPlugin_logic_machine_mie_mtie;
  reg                 PrivilegedPlugin_logic_machine_mie_msie;
  reg                 PrivilegedPlugin_logic_machine_medeleg_iam;
  reg                 PrivilegedPlugin_logic_machine_medeleg_bp;
  reg                 PrivilegedPlugin_logic_machine_medeleg_eu;
  reg                 PrivilegedPlugin_logic_machine_medeleg_es;
  reg                 PrivilegedPlugin_logic_machine_medeleg_ipf;
  reg                 PrivilegedPlugin_logic_machine_medeleg_lpf;
  reg                 PrivilegedPlugin_logic_machine_medeleg_spf;
  reg                 PrivilegedPlugin_logic_machine_mideleg_st;
  reg                 PrivilegedPlugin_logic_machine_mideleg_se;
  reg                 PrivilegedPlugin_logic_machine_mideleg_ss;
  reg                 PrivilegedPlugin_logic_supervisor_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_supervisor_cause_code;
  reg                 PrivilegedPlugin_logic_supervisor_sstatus_sie;
  reg                 PrivilegedPlugin_logic_supervisor_sstatus_spie;
  reg        [0:0]    PrivilegedPlugin_logic_supervisor_sstatus_spp;
  reg                 PrivilegedPlugin_logic_supervisor_sip_seipSoft;
  reg                 PrivilegedPlugin_logic_supervisor_sip_seipInput;
  wire                PrivilegedPlugin_logic_supervisor_sip_seipOr;
  reg                 PrivilegedPlugin_logic_supervisor_sip_stip;
  reg                 PrivilegedPlugin_logic_supervisor_sip_ssip;
  wire                PrivilegedPlugin_logic_supervisor_sip_seipMasked;
  wire                PrivilegedPlugin_logic_supervisor_sip_stipMasked;
  wire                PrivilegedPlugin_logic_supervisor_sip_ssipMasked;
  reg                 PrivilegedPlugin_logic_supervisor_sie_seie;
  reg                 PrivilegedPlugin_logic_supervisor_sie_stie;
  reg                 PrivilegedPlugin_logic_supervisor_sie_ssie;
  wire                _zz_when_PrivilegedPlugin_l637;
  wire                _zz_when_PrivilegedPlugin_l637_1;
  wire                _zz_when_PrivilegedPlugin_l637_2;
  reg                 PrivilegedPlugin_logic_rescheduleUnbuffered_valid;
  reg                 PrivilegedPlugin_logic_rescheduleUnbuffered_ready;
  reg        [3:0]    PrivilegedPlugin_logic_rescheduleUnbuffered_payload_cause;
  reg        [31:0]   PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc;
  reg        [31:0]   PrivilegedPlugin_logic_rescheduleUnbuffered_payload_tval;
  wire                PrivilegedPlugin_logic_rescheduleUnbuffered_payload_fromCommit;
  wire                PrivilegedPlugin_logic_reschedule_valid;
  reg                 PrivilegedPlugin_logic_reschedule_ready;
  wire       [3:0]    PrivilegedPlugin_logic_reschedule_payload_cause;
  wire       [31:0]   PrivilegedPlugin_logic_reschedule_payload_epc;
  wire       [31:0]   PrivilegedPlugin_logic_reschedule_payload_tval;
  wire                PrivilegedPlugin_logic_reschedule_payload_fromCommit;
  reg                 PrivilegedPlugin_logic_rescheduleUnbuffered_rValid;
  reg        [3:0]    PrivilegedPlugin_logic_rescheduleUnbuffered_rData_cause;
  reg        [31:0]   PrivilegedPlugin_logic_rescheduleUnbuffered_rData_epc;
  reg        [31:0]   PrivilegedPlugin_logic_rescheduleUnbuffered_rData_tval;
  reg                 PrivilegedPlugin_logic_rescheduleUnbuffered_rData_fromCommit;
  wire                when_Stream_l369;
  wire                when_PrivilegedPlugin_l585;
  wire                PrivilegedPlugin_logic_targetMachine;
  reg        [31:0]   PrivilegedPlugin_logic_readed;
  wire                PerformanceCounterPlugin_logic_branchMissEvent;
  reg                 _zz_PerformanceCounterPlugin_logic_branchMissEvent;
  reg        [1:0]    PerformanceCounterPlugin_logic_commitCount;
  reg                 PerformanceCounterPlugin_logic_ignoreNextCommit;
  wire                when_PerformanceCounterPlugin_l65;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_0;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_1;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_2;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_3;
  reg        [5:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded;
  reg        [5:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_1;
  reg        [5:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2;
  reg        [1:0]    PerformanceCounterPlugin_logic_commitCount_regNext;
  reg        [5:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3;
  reg        [5:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4;
  reg        [5:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5;
  reg        [5:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6;
  reg        [2:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_7;
  reg        [2:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_8;
  reg        [2:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_9;
  reg        [2:0]    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_10;
  wire                PerformanceCounterPlugin_logic_fsm_wantExit;
  reg                 PerformanceCounterPlugin_logic_fsm_wantStart;
  wire                PerformanceCounterPlugin_logic_fsm_wantKill;
  wire                PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid;
  reg                 PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready;
  wire       [2:0]    PerformanceCounterPlugin_logic_fsm_csrReadCmd_payload_address;
  wire                PerformanceCounterPlugin_logic_fsm_flusherCmd_valid;
  reg                 PerformanceCounterPlugin_logic_fsm_flusherCmd_ready;
  wire       [2:0]    PerformanceCounterPlugin_logic_fsm_flusherCmd_payload_address;
  reg                 PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid;
  reg                 PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready;
  wire       [2:0]    PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address;
  wire                PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_high;
  reg                 PerformanceCounterPlugin_logic_fsm_cmd_flusher;
  reg        [2:0]    PerformanceCounterPlugin_logic_fsm_cmd_address;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_valid;
  wire                ALU0_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   ALU0_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [2:0]    ALU0_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   ALU0_IntFormatPlugin_logic_stages_0_raw;
  reg        [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  reg        [31:0]   _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  reg        [31:0]   ALU0_SrcPlugin_logic_addsub_rs2Patched;
  reg        [31:0]   ALU0_IntAluPlugin_logic_process_bitwise;
  reg        [31:0]   ALU0_IntAluPlugin_logic_process_result;
  wire       [4:0]    ALU0_ShiftPlugin_logic_process_amplitude;
  wire       [31:0]   ALU0_ShiftPlugin_logic_process_reversed;
  wire       [31:0]   ALU0_ShiftPlugin_logic_process_shifted;
  wire       [31:0]   ALU0_ShiftPlugin_logic_process_patched;
  wire       [2:0]    switch_Misc_l232;
  reg                 _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
  reg                 _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1;
  reg        [31:0]   ALU0_BranchPlugin_logic_process_target_a;
  reg        [31:0]   ALU0_BranchPlugin_logic_process_target_b;
  wire       [1:0]    ALU0_BranchPlugin_logic_process_slices;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_2_valid;
  wire                EU0_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   EU0_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [2:0]    EU0_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   EU0_IntFormatPlugin_logic_stages_0_raw;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  reg        [31:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_valid;
  reg                 _zz_EU0_ExecutionUnitBase_pipeline_execute_1_valid;
  reg        [31:0]   EU0_SrcPlugin_logic_addsub_rs2Patched;
  wire                EU0_MulPlugin_logic_wake_wakeRobsSel;
  wire                EU0_MulPlugin_logic_wake_wakeRegFileSel;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_valid;
  reg                 _zz_EU0_ExecutionUnitBase_pipeline_execute_2_valid;
  reg        [60:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0;
  reg        [60:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_1;
  reg        [60:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_2;
  reg        [2:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1;
  reg        [2:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_1;
  reg        [2:0]    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_2;
  reg        [65:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0;
  reg        [65:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0_1;
  wire                EU0_DivPlugin_logic_wake_wakeRobsSel;
  wire                EU0_DivPlugin_logic_wake_wakeRegFileSel;
  reg                 EU0_DivPlugin_logic_feed_cmdSent;
  wire                toplevel_EU0_DivPlugin_logic_div_io_cmd_fire;
  wire                when_DivPlugin_l76;
  wire                EU0_ExecutionUnitBase_pipeline_execute_0_haltRequest_DivPlugin_l83;
  wire                EU0_ExecutionUnitBase_pipeline_execute_1_haltRequest_DivPlugin_l91;
  wire       [34:0]   EU0_DivPlugin_logic_rsp_selected;
  wire       [34:0]   _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT;
  wire       [2:0]    AguPlugin_logic_func3;
  reg                 AguPlugin_logic_fired;
  wire                when_AguPlugin_l89;
  wire       [1:0]    EnvCallPlugin_logic_xretPriv;
  wire                when_EnvCallPlugin_l95;
  wire                when_EnvCallPlugin_l108;
  wire                EnvCallPlugin_logic_flushes_wantExit;
  reg                 EnvCallPlugin_logic_flushes_wantStart;
  wire                EnvCallPlugin_logic_flushes_wantKill;
  wire                FetchPlugin_stages_0_haltRequest_EnvCallPlugin_l125;
  reg                 EnvCallPlugin_logic_flushes_vmaInv;
  reg                 EnvCallPlugin_logic_flushes_fetchInv;
  reg                 EnvCallPlugin_logic_flushes_flushData;
  reg        [2:0]    EnvCallPlugin_logic_flushes_stateReg;
  reg        [2:0]    EnvCallPlugin_logic_flushes_stateNext;
  wire                when_EnvCallPlugin_l135;
  wire                EU0_CsrAccessPlugin_logic_wake_wakeRobsSel;
  wire                EU0_CsrAccessPlugin_logic_wake_wakeRegFileSel;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_valid;
  wire                ALU1_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   ALU1_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [2:0]    ALU1_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   ALU1_IntFormatPlugin_logic_stages_0_raw;
  reg        [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  reg        [31:0]   _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  reg        [31:0]   ALU1_SrcPlugin_logic_addsub_rs2Patched;
  reg        [31:0]   ALU1_IntAluPlugin_logic_process_bitwise;
  reg        [31:0]   ALU1_IntAluPlugin_logic_process_result;
  wire       [4:0]    ALU1_ShiftPlugin_logic_process_amplitude;
  wire       [31:0]   ALU1_ShiftPlugin_logic_process_reversed;
  wire       [31:0]   ALU1_ShiftPlugin_logic_process_shifted;
  wire       [31:0]   ALU1_ShiftPlugin_logic_process_patched;
  wire       [2:0]    switch_Misc_l232_1;
  reg                 _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
  reg                 _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1;
  reg        [31:0]   ALU1_BranchPlugin_logic_process_target_a;
  reg        [31:0]   ALU1_BranchPlugin_logic_process_target_b;
  wire       [1:0]    ALU1_BranchPlugin_logic_process_slices;
  wire                FrontendPlugin_allocated_haltRequest_FrontendPlugin_l67;
  wire                integer_RfTranslationPlugin_logic_onCommit_writeRd_0;
  wire                integer_RfTranslationPlugin_logic_onCommit_writeRd_1;
  wire       [5:0]    integer_RfTranslationPlugin_logic_onCommit_physRd_0;
  wire       [5:0]    integer_RfTranslationPlugin_logic_onCommit_physRd_1;
  wire       [4:0]    integer_RfTranslationPlugin_logic_onCommit_archRd_0;
  wire       [4:0]    integer_RfTranslationPlugin_logic_onCommit_archRd_1;
  reg        [5:0]    integer_RfTranslationPlugin_logic_init_counter;
  wire                integer_RfTranslationPlugin_logic_init_busy;
  wire                when_RfTranslationPlugin_l193;
  wire                when_RfTranslationPlugin_l193_1;
  wire                _zz_when_RfTranslationPlugin_l214;
  wire                when_RfTranslationPlugin_l214;
  wire                when_RfTranslationPlugin_l218;
  wire                when_RfTranslationPlugin_l218_1;
  wire                integer_RfAllocationPlugin_logic_push_mask_0;
  wire                integer_RfAllocationPlugin_logic_push_mask_1;
  wire                integer_RfAllocationPlugin_logic_push_writeRd_0;
  wire                integer_RfAllocationPlugin_logic_push_writeRd_1;
  wire       [5:0]    integer_RfAllocationPlugin_logic_push_physicalRdNew_0;
  wire       [5:0]    integer_RfAllocationPlugin_logic_push_physicalRdNew_1;
  wire       [5:0]    integer_RfAllocationPlugin_logic_push_physicalRdOld_0;
  wire       [5:0]    integer_RfAllocationPlugin_logic_push_physicalRdOld_1;
  wire                when_RfAllocationPlugin_l81;
  wire                when_RfAllocationPlugin_l81_1;
  reg        [6:0]    integer_RfAllocationPlugin_logic_init_counter;
  wire                integer_RfAllocationPlugin_logic_init_busy;
  wire                BranchContextPlugin_logic_onCommit_isBranch_0;
  wire                BranchContextPlugin_logic_onCommit_isBranch_1;
  wire                BranchContextPlugin_logic_onCommit_isBranchCommit_0;
  wire                BranchContextPlugin_logic_onCommit_isBranchCommit_1;
  wire       [4:0]    BranchContextPlugin_logic_onCommit_commitedNext;
  wire                HistoryPlugin_logic_onCommit_isConditionalBranch_0;
  wire                HistoryPlugin_logic_onCommit_isConditionalBranch_1;
  wire                HistoryPlugin_logic_onCommit_isTaken_0;
  wire                HistoryPlugin_logic_onCommit_isTaken_1;
  wire       [23:0]   HistoryPlugin_logic_onCommit_valueNext;
  wire                when_HistoryPlugin_l90;
  wire                when_HistoryPlugin_l90_1;
  reg        [23:0]   HistoryPlugin_logic_onFetch_value;
  reg        [23:0]   HistoryPlugin_logic_onFetch_valueNext;
  wire       [23:0]   HistoryPlugin_logic_update_pushes_0_stateNext;
  wire                when_HistoryPlugin_l115;
  wire       [23:0]   HistoryPlugin_logic_update_pushes_2_stateNext;
  wire                when_HistoryPlugin_l115_1;
  wire                when_HistoryPlugin_l115_2;
  wire       [23:0]   HistoryPlugin_logic_update_rescheduleFlush_instHistory;
  wire                HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch;
  wire                HistoryPlugin_logic_update_rescheduleFlush_isTaken;
  wire       [23:0]   HistoryPlugin_logic_update_rescheduleFlush_newHistory;
  wire       [3:0]    DecoderPredictionPlugin_logic_ras_healPush;
  wire       [3:0]    DecoderPredictionPlugin_logic_ras_healPop;
  wire                DecoderPredictionPlugin_logic_decodePatch_rasPushUsed;
  wire                Lsu2Plugin_logic_translationWake;
  wire                Lsu2Plugin_logic_sqWritebackEvent_valid;
  wire       [3:0]    Lsu2Plugin_logic_sqWritebackEvent_payload;
  wire                Lsu2Plugin_logic_sqFeedEvent_valid;
  wire       [3:0]    Lsu2Plugin_logic_sqFeedEvent_payload;
  reg                 Lsu2Plugin_logic_lq_regs_0_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_0_valid;
  reg                 Lsu2Plugin_logic_lq_regs_0_redo;
  reg                 Lsu2Plugin_logic_lq_regs_0_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_0_delete;
  reg                 Lsu2Plugin_logic_lq_regs_0_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_0_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_0_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_0_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315;
  wire                when_Lsu2Plugin_l338;
  reg                 Lsu2Plugin_logic_lq_regs_1_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_1_valid;
  reg                 Lsu2Plugin_logic_lq_regs_1_redo;
  reg                 Lsu2Plugin_logic_lq_regs_1_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_1_delete;
  reg                 Lsu2Plugin_logic_lq_regs_1_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_1_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_1_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_1_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_1_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_1;
  wire                when_Lsu2Plugin_l338_1;
  reg                 Lsu2Plugin_logic_lq_regs_2_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_2_valid;
  reg                 Lsu2Plugin_logic_lq_regs_2_redo;
  reg                 Lsu2Plugin_logic_lq_regs_2_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_2_delete;
  reg                 Lsu2Plugin_logic_lq_regs_2_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_2_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_2_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_2_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_2_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_2;
  wire                when_Lsu2Plugin_l338_2;
  reg                 Lsu2Plugin_logic_lq_regs_3_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_3_valid;
  reg                 Lsu2Plugin_logic_lq_regs_3_redo;
  reg                 Lsu2Plugin_logic_lq_regs_3_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_3_delete;
  reg                 Lsu2Plugin_logic_lq_regs_3_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_3_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_3_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_3_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_3_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_3;
  wire                when_Lsu2Plugin_l338_3;
  reg                 Lsu2Plugin_logic_lq_regs_4_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_4_valid;
  reg                 Lsu2Plugin_logic_lq_regs_4_redo;
  reg                 Lsu2Plugin_logic_lq_regs_4_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_4_delete;
  reg                 Lsu2Plugin_logic_lq_regs_4_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_4_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_4_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_4_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_4_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_4;
  wire                when_Lsu2Plugin_l338_4;
  reg                 Lsu2Plugin_logic_lq_regs_5_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_5_valid;
  reg                 Lsu2Plugin_logic_lq_regs_5_redo;
  reg                 Lsu2Plugin_logic_lq_regs_5_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_5_delete;
  reg                 Lsu2Plugin_logic_lq_regs_5_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_5_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_5_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_5_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_5_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_5;
  wire                when_Lsu2Plugin_l338_5;
  reg                 Lsu2Plugin_logic_lq_regs_6_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_6_valid;
  reg                 Lsu2Plugin_logic_lq_regs_6_redo;
  reg                 Lsu2Plugin_logic_lq_regs_6_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_6_delete;
  reg                 Lsu2Plugin_logic_lq_regs_6_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_6_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_6_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_6_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_6_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_6;
  wire                when_Lsu2Plugin_l338_6;
  reg                 Lsu2Plugin_logic_lq_regs_7_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_7_valid;
  reg                 Lsu2Plugin_logic_lq_regs_7_redo;
  reg                 Lsu2Plugin_logic_lq_regs_7_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_7_delete;
  reg                 Lsu2Plugin_logic_lq_regs_7_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_7_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_7_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_7_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_7_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_7;
  wire                when_Lsu2Plugin_l338_7;
  reg                 Lsu2Plugin_logic_lq_regs_8_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_8_valid;
  reg                 Lsu2Plugin_logic_lq_regs_8_redo;
  reg                 Lsu2Plugin_logic_lq_regs_8_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_8_delete;
  reg                 Lsu2Plugin_logic_lq_regs_8_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_8_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_8_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_8_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_8_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_8_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_8_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_8;
  wire                when_Lsu2Plugin_l338_8;
  reg                 Lsu2Plugin_logic_lq_regs_9_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_9_valid;
  reg                 Lsu2Plugin_logic_lq_regs_9_redo;
  reg                 Lsu2Plugin_logic_lq_regs_9_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_9_delete;
  reg                 Lsu2Plugin_logic_lq_regs_9_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_9_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_9_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_9_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_9_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_9_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_9_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_9;
  wire                when_Lsu2Plugin_l338_9;
  reg                 Lsu2Plugin_logic_lq_regs_10_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_10_valid;
  reg                 Lsu2Plugin_logic_lq_regs_10_redo;
  reg                 Lsu2Plugin_logic_lq_regs_10_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_10_delete;
  reg                 Lsu2Plugin_logic_lq_regs_10_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_10_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_10_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_10_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_10_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_10_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_10_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_10;
  wire                when_Lsu2Plugin_l338_10;
  reg                 Lsu2Plugin_logic_lq_regs_11_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_11_valid;
  reg                 Lsu2Plugin_logic_lq_regs_11_redo;
  reg                 Lsu2Plugin_logic_lq_regs_11_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_11_delete;
  reg                 Lsu2Plugin_logic_lq_regs_11_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_11_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_11_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_11_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_11_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_11_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_11_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_11;
  wire                when_Lsu2Plugin_l338_11;
  reg                 Lsu2Plugin_logic_lq_regs_12_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_12_valid;
  reg                 Lsu2Plugin_logic_lq_regs_12_redo;
  reg                 Lsu2Plugin_logic_lq_regs_12_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_12_delete;
  reg                 Lsu2Plugin_logic_lq_regs_12_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_12_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_12_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_12_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_12_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_12_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_12_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_12;
  wire                when_Lsu2Plugin_l338_12;
  reg                 Lsu2Plugin_logic_lq_regs_13_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_13_valid;
  reg                 Lsu2Plugin_logic_lq_regs_13_redo;
  reg                 Lsu2Plugin_logic_lq_regs_13_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_13_delete;
  reg                 Lsu2Plugin_logic_lq_regs_13_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_13_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_13_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_13_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_13_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_13_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_13_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_13;
  wire                when_Lsu2Plugin_l338_13;
  reg                 Lsu2Plugin_logic_lq_regs_14_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_14_valid;
  reg                 Lsu2Plugin_logic_lq_regs_14_redo;
  reg                 Lsu2Plugin_logic_lq_regs_14_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_14_delete;
  reg                 Lsu2Plugin_logic_lq_regs_14_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_14_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_14_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_14_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_14_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_14_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_14_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_14;
  wire                when_Lsu2Plugin_l338_14;
  reg                 Lsu2Plugin_logic_lq_regs_15_allocation;
  reg                 Lsu2Plugin_logic_lq_regs_15_valid;
  reg                 Lsu2Plugin_logic_lq_regs_15_redo;
  reg                 Lsu2Plugin_logic_lq_regs_15_redoSet;
  reg                 Lsu2Plugin_logic_lq_regs_15_delete;
  reg                 Lsu2Plugin_logic_lq_regs_15_sqChecked;
  reg                 Lsu2Plugin_logic_lq_regs_15_niceHazard;
  reg        [9:0]    Lsu2Plugin_logic_lq_regs_15_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_15_address_mask;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefill;
  reg                 Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_lq_regs_15_waitOn_sqWriteback;
  reg                 Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeed;
  reg        [3:0]    Lsu2Plugin_logic_lq_regs_15_waitOn_sqId;
  reg        [1:0]    Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefillSet;
  reg                 Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAnySet;
  reg                 Lsu2Plugin_logic_lq_regs_15_waitOn_sqWritebackSet;
  reg                 Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeedSet;
  wire                when_Lsu2Plugin_l315_15;
  wire                when_Lsu2Plugin_l338_15;
  reg        [14:0]   Lsu2Plugin_logic_lq_ptr_priority;
  reg        [14:0]   Lsu2Plugin_logic_lq_ptr_priorityLast;
  reg        [4:0]    Lsu2Plugin_logic_lq_ptr_alloc;
  reg        [4:0]    Lsu2Plugin_logic_lq_ptr_free;
  wire       [3:0]    Lsu2Plugin_logic_lq_ptr_allocReal;
  wire       [3:0]    Lsu2Plugin_logic_lq_ptr_freeReal;
  reg        [4:0]    Lsu2Plugin_logic_lq_tracker_freeNext;
  reg        [4:0]    Lsu2Plugin_logic_lq_tracker_free;
  reg        [1:0]    _zz_Lsu2Plugin_logic_lq_tracker_freeReduced;
  wire                when_UInt_l120;
  reg        [1:0]    Lsu2Plugin_logic_lq_tracker_freeReduced;
  wire       [1:0]    Lsu2Plugin_logic_lq_tracker_add;
  reg        [1:0]    Lsu2Plugin_logic_lq_tracker_sub;
  reg                 Lsu2Plugin_logic_lq_tracker_clear;
  wire                Lsu2Plugin_logic_lq_onCommit_lqAlloc_0;
  wire                Lsu2Plugin_logic_lq_onCommit_lqAlloc_1;
  wire                Lsu2Plugin_logic_lq_onCommit_lqCommits_0;
  wire                Lsu2Plugin_logic_lq_onCommit_lqCommits_1;
  wire       [1:0]    Lsu2Plugin_logic_lq_onCommit_lqCommitCount;
  wire       [4:0]    Lsu2Plugin_logic_lq_onCommit_free;
  wire       [14:0]   Lsu2Plugin_logic_lq_onCommit_priority;
  wire                when_Lsu2Plugin_l454;
  wire                when_Lsu2Plugin_l454_1;
  wire                when_Lsu2Plugin_l454_2;
  wire                when_Lsu2Plugin_l454_3;
  wire                when_Lsu2Plugin_l454_4;
  wire                when_Lsu2Plugin_l454_5;
  wire                when_Lsu2Plugin_l454_6;
  wire                when_Lsu2Plugin_l454_7;
  wire                when_Lsu2Plugin_l454_8;
  wire                when_Lsu2Plugin_l454_9;
  wire                when_Lsu2Plugin_l454_10;
  wire                when_Lsu2Plugin_l454_11;
  wire                when_Lsu2Plugin_l454_12;
  wire                when_Lsu2Plugin_l454_13;
  wire                when_Lsu2Plugin_l454_14;
  wire                when_Lsu2Plugin_l454_15;
  wire                when_Lsu2Plugin_l454_16;
  wire                when_Lsu2Plugin_l454_17;
  wire                when_Lsu2Plugin_l454_18;
  wire                when_Lsu2Plugin_l454_19;
  wire                when_Lsu2Plugin_l454_20;
  wire                when_Lsu2Plugin_l454_21;
  wire                when_Lsu2Plugin_l454_22;
  wire                when_Lsu2Plugin_l454_23;
  wire                when_Lsu2Plugin_l454_24;
  wire                when_Lsu2Plugin_l454_25;
  wire                when_Lsu2Plugin_l454_26;
  wire                when_Lsu2Plugin_l454_27;
  wire                when_Lsu2Plugin_l454_28;
  wire                when_Lsu2Plugin_l454_29;
  wire                when_Lsu2Plugin_l454_30;
  wire                when_Lsu2Plugin_l454_31;
  reg                 Lsu2Plugin_logic_lq_reservation_kill;
  reg                 Lsu2Plugin_logic_lq_reservation_valid;
  reg        [31:0]   Lsu2Plugin_logic_lq_reservation_address;
  reg        [6:0]    Lsu2Plugin_logic_lq_reservation_counter;
  wire                when_Lsu2Plugin_l484;
  wire                Lsu2Plugin_logic_lq_hazardPrediction_hazard;
  reg                 Lsu2Plugin_logic_lq_hazardPrediction_write_valid;
  reg        [6:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address;
  reg        [2:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score;
  reg        [15:0]   Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag;
  reg        [3:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta;
  wire       [6:0]    _zz_when_MultiportRam_l362_2;
  wire       [22:0]   _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
  wire                Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_valid;
  wire       [6:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_address;
  wire       [2:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_score;
  wire       [15:0]   Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_tag;
  wire       [3:0]    Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_delta;
  wire                Lsu2Plugin_logic_lq_hitPrediction_hazard;
  wire                Lsu2Plugin_logic_lq_hitPrediction_write_valid;
  wire       [9:0]    Lsu2Plugin_logic_lq_hitPrediction_write_payload_address;
  wire       [5:0]    Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter;
  wire       [9:0]    _zz_when_MultiportRam_l362_3;
  wire       [5:0]    _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter;
  wire                Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_valid;
  wire       [9:0]    Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_address;
  wire       [5:0]    Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_data_counter;
  reg                 Lsu2Plugin_logic_sq_regs_0_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_0_valid;
  reg                 Lsu2Plugin_logic_sq_regs_0_redo;
  reg                 Lsu2Plugin_logic_sq_regs_0_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_0_delete;
  reg                 Lsu2Plugin_logic_sq_regs_0_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_0_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_0_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_0_commited;
  reg                 Lsu2Plugin_logic_sq_regs_0_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369;
  wire                when_Lsu2Plugin_l385;
  reg                 Lsu2Plugin_logic_sq_regs_1_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_1_valid;
  reg                 Lsu2Plugin_logic_sq_regs_1_redo;
  reg                 Lsu2Plugin_logic_sq_regs_1_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_1_delete;
  reg                 Lsu2Plugin_logic_sq_regs_1_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_1_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_1_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_1_commited;
  reg                 Lsu2Plugin_logic_sq_regs_1_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_1;
  wire                when_Lsu2Plugin_l385_1;
  reg                 Lsu2Plugin_logic_sq_regs_2_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_2_valid;
  reg                 Lsu2Plugin_logic_sq_regs_2_redo;
  reg                 Lsu2Plugin_logic_sq_regs_2_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_2_delete;
  reg                 Lsu2Plugin_logic_sq_regs_2_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_2_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_2_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_2_commited;
  reg                 Lsu2Plugin_logic_sq_regs_2_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_2;
  wire                when_Lsu2Plugin_l385_2;
  reg                 Lsu2Plugin_logic_sq_regs_3_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_3_valid;
  reg                 Lsu2Plugin_logic_sq_regs_3_redo;
  reg                 Lsu2Plugin_logic_sq_regs_3_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_3_delete;
  reg                 Lsu2Plugin_logic_sq_regs_3_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_3_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_3_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_3_commited;
  reg                 Lsu2Plugin_logic_sq_regs_3_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_3;
  wire                when_Lsu2Plugin_l385_3;
  reg                 Lsu2Plugin_logic_sq_regs_4_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_4_valid;
  reg                 Lsu2Plugin_logic_sq_regs_4_redo;
  reg                 Lsu2Plugin_logic_sq_regs_4_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_4_delete;
  reg                 Lsu2Plugin_logic_sq_regs_4_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_4_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_4_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_4_commited;
  reg                 Lsu2Plugin_logic_sq_regs_4_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_4;
  wire                when_Lsu2Plugin_l385_4;
  reg                 Lsu2Plugin_logic_sq_regs_5_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_5_valid;
  reg                 Lsu2Plugin_logic_sq_regs_5_redo;
  reg                 Lsu2Plugin_logic_sq_regs_5_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_5_delete;
  reg                 Lsu2Plugin_logic_sq_regs_5_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_5_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_5_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_5_commited;
  reg                 Lsu2Plugin_logic_sq_regs_5_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_5;
  wire                when_Lsu2Plugin_l385_5;
  reg                 Lsu2Plugin_logic_sq_regs_6_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_6_valid;
  reg                 Lsu2Plugin_logic_sq_regs_6_redo;
  reg                 Lsu2Plugin_logic_sq_regs_6_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_6_delete;
  reg                 Lsu2Plugin_logic_sq_regs_6_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_6_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_6_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_6_commited;
  reg                 Lsu2Plugin_logic_sq_regs_6_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_6;
  wire                when_Lsu2Plugin_l385_6;
  reg                 Lsu2Plugin_logic_sq_regs_7_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_7_valid;
  reg                 Lsu2Plugin_logic_sq_regs_7_redo;
  reg                 Lsu2Plugin_logic_sq_regs_7_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_7_delete;
  reg                 Lsu2Plugin_logic_sq_regs_7_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_7_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_7_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_7_commited;
  reg                 Lsu2Plugin_logic_sq_regs_7_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_7;
  wire                when_Lsu2Plugin_l385_7;
  reg                 Lsu2Plugin_logic_sq_regs_8_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_8_valid;
  reg                 Lsu2Plugin_logic_sq_regs_8_redo;
  reg                 Lsu2Plugin_logic_sq_regs_8_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_8_delete;
  reg                 Lsu2Plugin_logic_sq_regs_8_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_8_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_8_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_8_commited;
  reg                 Lsu2Plugin_logic_sq_regs_8_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_8;
  wire                when_Lsu2Plugin_l385_8;
  reg                 Lsu2Plugin_logic_sq_regs_9_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_9_valid;
  reg                 Lsu2Plugin_logic_sq_regs_9_redo;
  reg                 Lsu2Plugin_logic_sq_regs_9_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_9_delete;
  reg                 Lsu2Plugin_logic_sq_regs_9_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_9_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_9_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_9_commited;
  reg                 Lsu2Plugin_logic_sq_regs_9_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_9;
  wire                when_Lsu2Plugin_l385_9;
  reg                 Lsu2Plugin_logic_sq_regs_10_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_10_valid;
  reg                 Lsu2Plugin_logic_sq_regs_10_redo;
  reg                 Lsu2Plugin_logic_sq_regs_10_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_10_delete;
  reg                 Lsu2Plugin_logic_sq_regs_10_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_10_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_10_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_10_commited;
  reg                 Lsu2Plugin_logic_sq_regs_10_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_10;
  wire                when_Lsu2Plugin_l385_10;
  reg                 Lsu2Plugin_logic_sq_regs_11_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_11_valid;
  reg                 Lsu2Plugin_logic_sq_regs_11_redo;
  reg                 Lsu2Plugin_logic_sq_regs_11_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_11_delete;
  reg                 Lsu2Plugin_logic_sq_regs_11_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_11_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_11_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_11_commited;
  reg                 Lsu2Plugin_logic_sq_regs_11_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_11;
  wire                when_Lsu2Plugin_l385_11;
  reg                 Lsu2Plugin_logic_sq_regs_12_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_12_valid;
  reg                 Lsu2Plugin_logic_sq_regs_12_redo;
  reg                 Lsu2Plugin_logic_sq_regs_12_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_12_delete;
  reg                 Lsu2Plugin_logic_sq_regs_12_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_12_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_12_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_12_commited;
  reg                 Lsu2Plugin_logic_sq_regs_12_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_12;
  wire                when_Lsu2Plugin_l385_12;
  reg                 Lsu2Plugin_logic_sq_regs_13_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_13_valid;
  reg                 Lsu2Plugin_logic_sq_regs_13_redo;
  reg                 Lsu2Plugin_logic_sq_regs_13_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_13_delete;
  reg                 Lsu2Plugin_logic_sq_regs_13_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_13_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_13_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_13_commited;
  reg                 Lsu2Plugin_logic_sq_regs_13_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_13;
  wire                when_Lsu2Plugin_l385_13;
  reg                 Lsu2Plugin_logic_sq_regs_14_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_14_valid;
  reg                 Lsu2Plugin_logic_sq_regs_14_redo;
  reg                 Lsu2Plugin_logic_sq_regs_14_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_14_delete;
  reg                 Lsu2Plugin_logic_sq_regs_14_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_14_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_14_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_14_commited;
  reg                 Lsu2Plugin_logic_sq_regs_14_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_14;
  wire                when_Lsu2Plugin_l385_14;
  reg                 Lsu2Plugin_logic_sq_regs_15_allocation;
  reg                 Lsu2Plugin_logic_sq_regs_15_valid;
  reg                 Lsu2Plugin_logic_sq_regs_15_redo;
  reg                 Lsu2Plugin_logic_sq_regs_15_redoSet;
  reg                 Lsu2Plugin_logic_sq_regs_15_delete;
  reg                 Lsu2Plugin_logic_sq_regs_15_dataValid;
  reg        [9:0]    Lsu2Plugin_logic_sq_regs_15_address_pageOffset;
  reg        [3:0]    Lsu2Plugin_logic_sq_regs_15_address_mask;
  reg                 Lsu2Plugin_logic_sq_regs_15_commited;
  reg                 Lsu2Plugin_logic_sq_regs_15_commitedNext;
  reg                 Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAny;
  reg                 Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAnySet;
  wire                when_Lsu2Plugin_l369_15;
  wire                when_Lsu2Plugin_l385_15;
  reg                 Lsu2Plugin_logic_sq_mem_swap;
  reg        [2:0]    Lsu2Plugin_logic_sq_mem_op;
  reg        [5:0]    Lsu2Plugin_logic_sq_mem_physRd;
  reg                 Lsu2Plugin_logic_sq_mem_writeRd;
  reg        [14:0]   Lsu2Plugin_logic_sq_ptr_priority;
  reg        [14:0]   Lsu2Plugin_logic_sq_ptr_priorityLast;
  reg        [4:0]    Lsu2Plugin_logic_sq_ptr_alloc;
  reg        [4:0]    Lsu2Plugin_logic_sq_ptr_commit;
  reg        [4:0]    Lsu2Plugin_logic_sq_ptr_writeBack;
  reg        [4:0]    Lsu2Plugin_logic_sq_ptr_free;
  wire       [3:0]    Lsu2Plugin_logic_sq_ptr_allocReal;
  wire       [3:0]    Lsu2Plugin_logic_sq_ptr_freeReal /* verilator public */ ;
  wire       [3:0]    Lsu2Plugin_logic_sq_ptr_writeBackReal;
  wire       [3:0]    Lsu2Plugin_logic_sq_ptr_commitReal;
  wire       [4:0]    Lsu2Plugin_logic_sq_ptr_commitNext;
  reg                 Lsu2Plugin_logic_sq_ptr_onFree_valid;
  wire       [3:0]    Lsu2Plugin_logic_sq_ptr_onFree_payload;
  reg                 Lsu2Plugin_logic_sq_ptr_onFreeLast_valid;
  reg        [3:0]    Lsu2Plugin_logic_sq_ptr_onFreeLast_payload;
  wire                when_Lsu2Plugin_l572;
  wire       [4:0]    Lsu2Plugin_logic_sq_tracker_freeNext;
  reg        [4:0]    Lsu2Plugin_logic_sq_tracker_free;
  reg        [1:0]    _zz_Lsu2Plugin_logic_sq_tracker_freeReduced;
  wire                when_UInt_l120_1;
  reg        [1:0]    Lsu2Plugin_logic_sq_tracker_freeReduced;
  reg        [0:0]    Lsu2Plugin_logic_sq_tracker_add;
  reg        [1:0]    Lsu2Plugin_logic_sq_tracker_sub;
  wire                Lsu2Plugin_logic_sq_onCommit_sqAlloc_0;
  wire                Lsu2Plugin_logic_sq_onCommit_sqAlloc_1;
  wire       [0:0]    Lsu2Plugin_logic_sq_onCommit_sqCommits_0;
  wire       [0:0]    Lsu2Plugin_logic_sq_onCommit_sqCommits_1;
  wire       [4:0]    Lsu2Plugin_logic_sq_onCommit_commitComb;
  wire                when_Lsu2Plugin_l591;
  wire       [15:0]   _zz_45;
  wire                when_Lsu2Plugin_l591_1;
  wire       [15:0]   _zz_46;
  wire                Lsu2Plugin_logic_allocation_loads_requests_0;
  wire                Lsu2Plugin_logic_allocation_loads_requests_1;
  wire       [1:0]    Lsu2Plugin_logic_allocation_loads_requestsCount;
  wire                Lsu2Plugin_logic_allocation_loads_full;
  wire       [4:0]    Lsu2Plugin_logic_allocation_loads_alloc;
  wire                Lsu2Plugin_logic_allocation_stores_requests_0;
  wire                Lsu2Plugin_logic_allocation_stores_requests_1;
  wire       [1:0]    Lsu2Plugin_logic_allocation_stores_requestsCount;
  wire                Lsu2Plugin_logic_allocation_stores_full;
  wire       [4:0]    Lsu2Plugin_logic_allocation_stores_alloc;
  wire                FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l620;
  wire                FrontendPlugin_dispatch_isFireing /* verilator public */ ;
  wire                Lsu2Plugin_logic_aguPush_0_pushLq;
  wire                Lsu2Plugin_logic_aguPush_0_pushSq;
  reg        [3:0]    _zz_Lsu2Plugin_logic_aguPush_0_dataMask;
  wire       [3:0]    Lsu2Plugin_logic_aguPush_0_dataMask;
  wire       [3:0]    switch_Utils_l1437;
  wire                Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_valid;
  wire       [6:0]    Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_payload;
  wire       [2:0]    Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
  wire       [15:0]   Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_tag;
  wire       [3:0]    Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_delta;
  wire       [22:0]   _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_1;
  wire       [15:0]   Lsu2Plugin_logic_aguPush_0_hazardPrediction_hash;
  wire                Lsu2Plugin_logic_aguPush_0_hazardPrediction_hit;
  wire                Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_valid;
  wire       [9:0]    Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_payload;
  wire       [5:0]    Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter;
  wire                Lsu2Plugin_logic_aguPush_0_hitPrediction_likelyToHit;
  wire                when_Lsu2Plugin_l733;
  wire       [3:0]    switch_Utils_l1437_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_valid;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_input;
  wire       [14:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_priorityBits;
  wire       [30:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask;
  wire       [30:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_2;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_8;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_13;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_14;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_15;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_16;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_17;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_18;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_19;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_20;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_21;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_22;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_23;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_24;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_25;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_26;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_27;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_28;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_29;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_30;
  reg        [30:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_4;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_8;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_8;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_9_to_10;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_9_to_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_13;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_14;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_14;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_15_to_16;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_15_to_17;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_19;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_20;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_21_to_22;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_21_to_23;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_23;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_24_to_25;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_24_to_26;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_26;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_27_to_28;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_27_to_29;
  wire       [30:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pLow;
  wire       [14:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pHigh;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_input;
  wire       [14:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_priorityBits;
  wire       [30:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask;
  wire       [30:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_2;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_8;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_13;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_14;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_15;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_16;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_17;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_18;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_19;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_20;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_21;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_22;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_23;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_24;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_25;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_26;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_27;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_28;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_29;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_30;
  reg        [30:0]   _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_4;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_5;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_7;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_8;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_8;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_9_to_10;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_9_to_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_11;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_13;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_14;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_14;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_15_to_16;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_15_to_17;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_19;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_20;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_21_to_22;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_21_to_23;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_23;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_24_to_25;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_24_to_26;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_26;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_27_to_28;
  wire                Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_27_to_29;
  wire       [30:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pLow;
  wire       [14:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pHigh;
  wire       [15:0]   Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_1;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_3;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_7;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_8;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_9;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_10;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_11;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_12;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_13;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_14;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_15;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_16;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_17;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_18;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_1;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_3;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_7;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_8;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_9;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_10;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_11;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_12;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_13;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_14;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_15;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_16;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_17;
  wire                _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_18;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s1_valid;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_cmp;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_valid;
  reg                 _zz_Lsu2Plugin_logic_sharedPip_stages_1_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_1_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_2_valid;
  reg                 Lsu2Plugin_logic_sharedPip_stages_3_valid;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_wake;
  reg                 Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap;
  reg                 Lsu2Plugin_logic_sharedPip_speculateHitTrapRecovered;
  reg                 Lsu2Plugin_logic_sharedPip_speculativeHitPredictionGotReschedule;
  reg                 Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled;
  reg                 Lsu2Plugin_logic_sharedPip_feed_takeAgu;
  wire                when_Lsu2Plugin_l830;
  wire                when_Lsu2Plugin_l831;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l834;
  reg                 Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask;
  reg                 Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask;
  wire                when_Lsu2Plugin_l838;
  wire                when_Lsu2Plugin_l839;
  wire                when_Lsu2Plugin_l841;
  wire                Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842;
  wire                when_Lsu2Plugin_l843;
  wire                when_Lsu2Plugin_l845;
  wire                when_Lsu2Plugin_l849;
  wire                when_Lsu2Plugin_l920;
  wire                when_Lsu2Plugin_l929;
  wire       [3:0]    switch_Utils_l1437_2;
  wire       [3:0]    switch_Utils_l1437_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_isFireing;
  reg        [3:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT;
  wire                when_Lsu2Plugin_l959;
  wire                Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_valid;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_payload_robId;
  wire                Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_valid;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_payload_physical;
  wire                Lsu2Plugin_logic_sharedPip_stages_0_haltRequest_Lsu2Plugin_l990;
  wire                when_Lsu2Plugin_l997;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_loopback;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_youngerMask;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_olderMaskEmpty;
  reg        [15:0]   Lsu2Plugin_logic_sharedPip_checkSqMask_hits;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_8_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_8_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_9_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_9_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_10_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_10_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_11_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_11_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_12_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_12_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_13_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_13_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_14_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_14_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_15_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_entries_15_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkSqMask_olderHit;
  wire       [15:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input;
  wire       [14:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits;
  wire       [30:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask;
  wire       [30:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_1;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_2;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_8;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_13;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_14;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_15;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_16;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_17;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_18;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_19;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_20;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_21;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_22;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_23;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_24;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_25;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_26;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_27;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_28;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_29;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_30;
  reg        [30:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_4;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_10;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_16;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_17;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_19;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_22;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_25;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_26;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_28;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_29;
  wire       [30:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pLow;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pHigh;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_4;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_5;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_6;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_7;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_8;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_9;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_10;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_11;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_12;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_13;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_14;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel;
  wire                Lsu2Plugin_logic_sharedPip_stages_1_isFireing;
  wire                when_Lsu2Plugin_l1046;
  wire                when_Lsu2Plugin_l1052;
  wire                Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_addressMatch;
  wire                Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_fullMatch;
  wire                Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_translationFailure;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_data;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_checkLqHits_endId;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_checkLqHits_startMask;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_checkLqHits_endMask;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_loopback;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMaskEmpty;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_hit;
  wire                when_Lsu2Plugin_l1104;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_hit;
  wire                when_Lsu2Plugin_l1104_1;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_hit;
  wire                when_Lsu2Plugin_l1104_2;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_hit;
  wire                when_Lsu2Plugin_l1104_3;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_hit;
  wire                when_Lsu2Plugin_l1104_4;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_hit;
  wire                when_Lsu2Plugin_l1104_5;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_hit;
  wire                when_Lsu2Plugin_l1104_6;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_hit;
  wire                when_Lsu2Plugin_l1104_7;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_hit;
  wire                when_Lsu2Plugin_l1104_8;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_hit;
  wire                when_Lsu2Plugin_l1104_9;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_hit;
  wire                when_Lsu2Plugin_l1104_10;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_hit;
  wire                when_Lsu2Plugin_l1104_11;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_hit;
  wire                when_Lsu2Plugin_l1104_12;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_hit;
  wire                when_Lsu2Plugin_l1104_13;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_hit;
  wire                when_Lsu2Plugin_l1104_14;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_pageHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_wordHit;
  wire                Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_hit;
  wire                when_Lsu2Plugin_l1104_15;
  wire                Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerHit;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_input;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_priorityBits;
  wire       [30:0]   Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask;
  wire       [30:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_1;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_2;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_8;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_13;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_14;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_15;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_16;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_17;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_18;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_19;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_20;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_21;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_22;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_23;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_24;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_25;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_26;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_27;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_28;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_29;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_30;
  reg        [30:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_4;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_10;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_16;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_17;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_19;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_22;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_25;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_26;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_28;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_29;
  wire       [30:0]   Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pLow;
  wire       [14:0]   Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pHigh;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_4;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_5;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_6;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_7;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_8;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_9;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_10;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_11;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_12;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_13;
  wire                _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_14;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel;
  reg                 Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride;
  reg        [1:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress;
  reg                 Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_0;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_1;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_2;
  wire       [7:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted;
  wire                when_Lsu2Plugin_l1158;
  wire                _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
  reg        [31:0]   _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
  reg        [31:0]   _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3;
  wire       [31:0]   _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_4;
  reg        [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
  wire                Lsu2Plugin_logic_sharedPip_stages_2_isFireing;
  wire                Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_valid /* verilator public */ ;
  wire                Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_isLoad /* verilator public */ ;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_address /* verilator public */ ;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_readData /* verilator public */ ;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_robId /* verilator public */ ;
  wire       [3:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_lqId /* verilator public */ ;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_size /* verilator public */ ;
  wire                Lsu2Plugin_logic_sharedPip_cacheRsp_doIt;
  reg                 Lsu2Plugin_logic_sharedPip_cacheRsp_success;
  wire                when_Lsu2Plugin_l1203;
  wire                when_Lsu2Plugin_l1205;
  wire                when_Lsu2Plugin_l1207;
  wire                when_Lsu2Plugin_l1209;
  wire                when_Lsu2Plugin_l1211;
  wire                when_Lsu2Plugin_l1213;
  wire       [3:0]    _zz_Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC;
  reg                 Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_valid;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_payload_robId;
  reg                 Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid;
  reg        [5:0]    Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_payload_physical;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_ctrl_lqMask;
  wire       [15:0]   Lsu2Plugin_logic_sharedPip_ctrl_sqMask;
  reg                 Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire                _zz_133;
  wire                _zz_134;
  wire       [1:0]    Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
  wire                Lsu2Plugin_logic_sharedPip_ctrl_doCompletion;
  wire                Lsu2Plugin_logic_sharedPip_stages_3_isFireing;
  wire                when_Lsu2Plugin_l1313;
  wire       [3:0]    _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
  wire                when_Lsu2Plugin_l1314;
  wire                when_Lsu2Plugin_l1333;
  wire                when_Lsu2Plugin_l1335;
  wire                _zz_when_Lsu2Plugin_l1348;
  reg        [2:0]    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score;
  wire                when_Lsu2Plugin_l1348;
  wire                when_Lsu2Plugin_l1351;
  wire                when_Lsu2Plugin_l1374;
  wire       [5:0]    _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next;
  wire       [6:0]    Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next;
  reg        [5:0]    _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter;
  wire                when_SInt_l131;
  wire                when_SInt_l132;
  wire                when_SInt_l138;
  reg                 Lsu2Plugin_logic_writeback_generation;
  reg        [1:0]    Lsu2Plugin_logic_writeback_waitOn_refillSlot;
  reg                 Lsu2Plugin_logic_writeback_waitOn_refillSlotAny;
  wire                Lsu2Plugin_logic_writeback_waitOn_ready;
  reg        [1:0]    Lsu2Plugin_logic_writeback_waitOn_refillSlotSet;
  reg                 Lsu2Plugin_logic_writeback_waitOn_refillSlotAnySet;
  wire                Lsu2Plugin_logic_writeback_feed_holdPrefetch;
  wire                toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_valid;
  wire                toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready;
  wire       [31:0]   toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_payload;
  reg                 toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rValid;
  reg        [31:0]   toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rData;
  wire                when_Stream_l369_1;
  wire                _zz_toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready;
  wire                Lsu2Plugin_logic_writeback_feed_prediction_valid;
  wire       [31:0]   Lsu2Plugin_logic_writeback_feed_prediction_payload;
  wire                Lsu2Plugin_logic_writeback_feed_io;
  wire       [1:0]    Lsu2Plugin_logic_writeback_feed_size;
  reg        [31:0]   Lsu2Plugin_logic_writeback_feed_data;
  reg                 Lsu2Plugin_logic_writeback_feed_skip;
  wire                Lsu2Plugin_logic_writeback_feed_doit;
  reg                 Lsu2Plugin_logic_writeback_feed_fire;
  reg        [3:0]    _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_valid;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_fault;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlot;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_generationKo;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_flush;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_prefetch;
  wire       [31:0]   Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_address;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_io;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_valid;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_fault;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlot;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_generationKo;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_flush;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_prefetch;
  wire       [31:0]   Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_address;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_io;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_valid;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_fault;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_redo;
  wire       [1:0]    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlot;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlotAny;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_generationKo;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_flush;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_prefetch;
  wire       [31:0]   Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_address;
  wire                Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_io;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_valid;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_fault;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_redo;
  reg        [1:0]    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlot;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlotAny;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_generationKo;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_flush;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_prefetch;
  reg        [31:0]   Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_address;
  reg                 Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_io;
  reg                 Lsu2Plugin_logic_writeback_rsp_whitebox_valid /* verilator public */ ;
  wire                when_Lsu2Plugin_l1488;
  wire                when_Lsu2Plugin_l1498;
  wire                when_Lsu2Plugin_l1509;
  wire                when_Lsu2Plugin_l1521;
  wire                when_Lsu2Plugin_l1524;
  wire                when_Lsu2Plugin_l1524_1;
  wire                when_Lsu2Plugin_l1524_2;
  wire                when_Lsu2Plugin_l1524_3;
  wire                when_Lsu2Plugin_l1524_4;
  wire                when_Lsu2Plugin_l1524_5;
  wire                when_Lsu2Plugin_l1524_6;
  wire                when_Lsu2Plugin_l1524_7;
  wire                when_Lsu2Plugin_l1524_8;
  wire                when_Lsu2Plugin_l1524_9;
  wire                when_Lsu2Plugin_l1524_10;
  wire                when_Lsu2Plugin_l1524_11;
  wire                when_Lsu2Plugin_l1524_12;
  wire                when_Lsu2Plugin_l1524_13;
  wire                when_Lsu2Plugin_l1524_14;
  wire                when_Lsu2Plugin_l1524_15;
  reg                 Lsu2Plugin_logic_flush_busy;
  reg                 Lsu2Plugin_logic_flush_doit;
  reg                 Lsu2Plugin_logic_flush_withFree;
  reg        [6:0]    Lsu2Plugin_logic_flush_cmdPtr;
  reg        [6:0]    Lsu2Plugin_logic_flush_rspPtr;
  wire                FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548;
  wire                when_Lsu2Plugin_l1553;
  wire                Lsu2Plugin_setup_cacheStore_cmd_fire;
  wire                when_Lsu2Plugin_l1561;
  wire                when_Lsu2Plugin_l1569;
  wire                Lsu2Plugin_logic_special_lqOnTop;
  wire                Lsu2Plugin_logic_special_sqOnTop;
  wire                Lsu2Plugin_logic_special_storeWriteBackUsable;
  wire                Lsu2Plugin_logic_special_storeSpecial;
  wire                Lsu2Plugin_logic_special_loadSpecial;
  wire                Lsu2Plugin_logic_special_storeHit;
  wire                Lsu2Plugin_logic_special_loadHit;
  wire                Lsu2Plugin_logic_special_hit;
  reg                 LsuPlugin_peripheralBus_rsp_valid_regNext;
  reg                 Lsu2Plugin_logic_special_fire;
  reg                 Lsu2Plugin_logic_special_enabled;
  reg                 Lsu2Plugin_logic_special_isStore;
  reg                 Lsu2Plugin_logic_special_isLoad;
  reg                 Lsu2Plugin_logic_special_cmdSent;
  wire                LsuPlugin_peripheralBus_cmd_fire;
  reg        [5:0]    Lsu2Plugin_logic_special_robId /* verilator public */ ;
  reg        [5:0]    Lsu2Plugin_logic_special_loadPhysRd;
  reg        [31:0]   Lsu2Plugin_logic_special_loadAddress;
  reg        [31:0]   Lsu2Plugin_logic_special_loadAddressVirt;
  reg        [1:0]    Lsu2Plugin_logic_special_loadSize;
  reg                 Lsu2Plugin_logic_special_loadUnsigned;
  reg                 Lsu2Plugin_logic_special_loadWriteRd;
  reg        [31:0]   Lsu2Plugin_logic_special_storeAddress;
  reg        [31:0]   Lsu2Plugin_logic_special_storeAddressVirt;
  reg        [1:0]    Lsu2Plugin_logic_special_storeSize;
  reg        [31:0]   Lsu2Plugin_logic_special_storeData;
  reg        [3:0]    Lsu2Plugin_logic_special_storeMask;
  reg                 Lsu2Plugin_logic_special_storeAmo;
  reg                 Lsu2Plugin_logic_special_storeSc;
  wire       [31:0]   Lsu2Plugin_logic_special_address;
  wire       [31:0]   Lsu2Plugin_logic_special_addressVirt;
  wire                Lsu2Plugin_logic_special_isIo;
  wire                Lsu2Plugin_logic_special_isAtomic;
  reg                 Lsu2Plugin_logic_special_wakeRob_valid;
  wire       [5:0]    Lsu2Plugin_logic_special_wakeRob_payload_robId;
  reg                 Lsu2Plugin_logic_special_wakeRf_valid;
  wire       [5:0]    Lsu2Plugin_logic_special_wakeRf_payload_physical;
  wire                Lsu2Plugin_logic_special_atomic_wantExit;
  reg                 Lsu2Plugin_logic_special_atomic_wantStart;
  wire                Lsu2Plugin_logic_special_atomic_wantKill;
  reg        [31:0]   Lsu2Plugin_logic_special_atomic_readed;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub;
  wire       [31:0]   _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1;
  wire                Lsu2Plugin_logic_special_atomic_alu_compare;
  wire                Lsu2Plugin_logic_special_atomic_alu_unsigned;
  wire       [31:0]   Lsu2Plugin_logic_special_atomic_alu_addSub;
  wire                Lsu2Plugin_logic_special_atomic_alu_less;
  wire                Lsu2Plugin_logic_special_atomic_alu_selectRf;
  wire       [2:0]    switch_Misc_l232_2;
  reg        [31:0]   Lsu2Plugin_logic_special_atomic_alu_raw;
  wire       [31:0]   Lsu2Plugin_logic_special_atomic_alu_result /* verilator public */ ;
  reg        [31:0]   Lsu2Plugin_logic_special_atomic_result;
  wire                when_Lsu2Plugin_l1683;
  wire                when_Lsu2Plugin_l1698;
  reg                 Lsu2Plugin_logic_special_atomic_gotReservation;
  reg        [1:0]    Lsu2Plugin_logic_special_atomic_lockDelayCounter;
  reg                 Lsu2Plugin_logic_special_atomic_comp_wakeRf;
  reg                 Lsu2Plugin_logic_special_atomic_comp_rfWrite;
  reg                 Lsu2Plugin_logic_special_atomic_loadWhitebox_valid /* verilator public */ ;
  wire       [31:0]   Lsu2Plugin_logic_special_atomic_loadWhitebox_readData /* verilator public */ ;
  reg                 Lsu2Plugin_logic_special_atomic_storeWhitebox_valid /* verilator public */ ;
  wire                Lsu2Plugin_logic_special_atomic_storeWhitebox_isSc /* verilator public */ ;
  wire                Lsu2Plugin_logic_special_atomic_storeWhitebox_scPassed /* verilator public */ ;
  wire                FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l1834;
  reg                 Lsu2Plugin_logic_lqFlush /* verilator public */ ;
  wire                when_Lsu2Plugin_l1909;
  wire                when_Lsu2Plugin_l1909_1;
  wire                when_Lsu2Plugin_l1909_2;
  wire                when_Lsu2Plugin_l1909_3;
  wire                when_Lsu2Plugin_l1909_4;
  wire                when_Lsu2Plugin_l1909_5;
  wire                when_Lsu2Plugin_l1909_6;
  wire                when_Lsu2Plugin_l1909_7;
  wire                when_Lsu2Plugin_l1909_8;
  wire                when_Lsu2Plugin_l1909_9;
  wire                when_Lsu2Plugin_l1909_10;
  wire                when_Lsu2Plugin_l1909_11;
  wire                when_Lsu2Plugin_l1909_12;
  wire                when_Lsu2Plugin_l1909_13;
  wire                when_Lsu2Plugin_l1909_14;
  wire                when_Lsu2Plugin_l1909_15;
  wire                sqAlloc_0_valid /* verilator public */ ;
  wire       [3:0]    sqAlloc_0_id /* verilator public */ ;
  wire                sqAlloc_1_valid /* verilator public */ ;
  wire       [3:0]    sqAlloc_1_id /* verilator public */ ;
  wire                sqFree_valid /* verilator public */ ;
  wire       [3:0]    sqFree_payload /* verilator public */ ;
  wire       [32:0]   _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken;
  reg                 ALU0_ExecutionUnitBase_pipeline_execute_1_valid;
  wire                ALU0_BranchPlugin_logic_branch_badEarlyTaken;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_1_isFireing;
  wire                ALU0_BranchPlugin_logic_branch_finalBranch_valid;
  wire       [3:0]    ALU0_BranchPlugin_logic_branch_finalBranch_payload_address;
  wire       [31:0]   ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice;
  wire       [31:0]   ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcTarget;
  wire                ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_taken;
  wire       [32:0]   _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken;
  reg                 ALU1_ExecutionUnitBase_pipeline_execute_1_valid;
  wire                ALU1_BranchPlugin_logic_branch_badEarlyTaken;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_1_isFireing;
  wire                ALU1_BranchPlugin_logic_branch_finalBranch_valid;
  wire       [3:0]    ALU1_BranchPlugin_logic_branch_finalBranch_payload_address;
  wire       [31:0]   ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice;
  wire       [31:0]   ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcTarget;
  wire                ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_taken;
  reg        [0:0]    MmuPlugin_logic_satp_mode;
  reg        [19:0]   MmuPlugin_logic_satp_ppn;
  reg                 MmuPlugin_logic_status_mxr;
  reg                 MmuPlugin_logic_status_sum;
  reg                 MmuPlugin_logic_status_mprv;
  wire       [0:0]    MmuPlugin_logic_satpModeWrite;
  reg                 FetchCachePlugin_setup_translationStorage_logic_refillOngoing;
  reg        [3:0]    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask;
  reg        [4:0]    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault;
  reg        [14:0]   FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willClear;
  reg        [1:0]    FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [1:0]    FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [1:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask;
  reg        [4:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault;
  reg        [4:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [9:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willClear;
  reg        [0:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_valueNext;
  reg        [0:0]    FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflow;
  reg                 Lsu2Plugin_setup_translationStorage_logic_refillOngoing;
  reg        [3:0]    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask;
  reg        [4:0]    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault;
  reg        [14:0]   Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willClear;
  reg        [1:0]    Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [1:0]    Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [1:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask;
  reg        [4:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault;
  reg        [4:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [9:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willClear;
  reg        [0:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_valueNext;
  reg        [0:0]    Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflow;
  reg                 Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg;
  wire                when_MmuPlugin_l260;
  reg                 Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg;
  wire                when_MmuPlugin_l260_1;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress;
  wire       [41:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid;
  wire       [41:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid;
  wire       [41:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid;
  wire       [41:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid;
  wire       [4:0]    Lsu2Plugin_logic_sharedPip_translationPort_logic_read_1_readAddress;
  wire       [21:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid;
  wire       [21:0]   _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hit;
  wire       [5:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_3;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_4;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_5;
  reg        [5:0]    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_1;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_2;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_3;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_4;
  wire       [5:0]    Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4;
  wire                _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException;
  wire       [31:0]   Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault;
  reg                 Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_needRefill;
  wire                Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_askRefill;
  wire                when_MmuPlugin_l297;
  wire                when_MmuPlugin_l298;
  wire                when_MmuPlugin_l300;
  wire                CsrRamPlugin_setup_initPort_valid;
  wire                CsrRamPlugin_setup_initPort_ready;
  wire       [4:0]    CsrRamPlugin_setup_initPort_address;
  wire       [31:0]   CsrRamPlugin_setup_initPort_data;
  reg                 PrivilegedPlugin_setup_ramRead_valid;
  wire                PrivilegedPlugin_setup_ramRead_ready;
  reg        [4:0]    PrivilegedPlugin_setup_ramRead_address;
  wire       [31:0]   PrivilegedPlugin_setup_ramRead_data;
  reg                 PrivilegedPlugin_setup_ramWrite_valid;
  wire                PrivilegedPlugin_setup_ramWrite_ready;
  reg        [4:0]    PrivilegedPlugin_setup_ramWrite_address;
  reg        [31:0]   PrivilegedPlugin_setup_ramWrite_data;
  reg                 PerformanceCounterPlugin_setup_readPort_valid;
  wire                PerformanceCounterPlugin_setup_readPort_ready;
  reg        [4:0]    PerformanceCounterPlugin_setup_readPort_address;
  wire       [31:0]   PerformanceCounterPlugin_setup_readPort_data;
  reg                 PerformanceCounterPlugin_setup_writePort_valid;
  wire                PerformanceCounterPlugin_setup_writePort_ready;
  reg        [4:0]    PerformanceCounterPlugin_setup_writePort_address;
  reg        [31:0]   PerformanceCounterPlugin_setup_writePort_data;
  reg                 PrivilegedPlugin_logic_interrupt_valid;
  reg        [3:0]    PrivilegedPlugin_logic_interrupt_code;
  reg        [1:0]    PrivilegedPlugin_logic_interrupt_targetPrivilege;
  wire                when_PrivilegedPlugin_l631;
  wire                when_PrivilegedPlugin_l631_1;
  wire                when_PrivilegedPlugin_l637;
  wire                when_PrivilegedPlugin_l637_1;
  wire                when_PrivilegedPlugin_l637_2;
  wire                when_PrivilegedPlugin_l637_3;
  wire                when_PrivilegedPlugin_l637_4;
  wire                when_PrivilegedPlugin_l637_5;
  wire                when_PrivilegedPlugin_l637_6;
  wire                when_PrivilegedPlugin_l637_7;
  wire                when_PrivilegedPlugin_l637_8;
  reg                 PrivilegedPlugin_logic_decoderInterrupt_raised;
  reg                 PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt;
  reg        [2:0]    PrivilegedPlugin_logic_decoderInterrupt_counter;
  wire                PrivilegedPlugin_logic_decoderInterrupt_doIt;
  wire                when_PrivilegedPlugin_l668;
  wire                when_PrivilegedPlugin_l672;
  wire                PrivilegedPlugin_logic_decoderInterrupt_buffer_sample;
  reg        [3:0]    PrivilegedPlugin_logic_decoderInterrupt_buffer_code;
  reg        [1:0]    PrivilegedPlugin_logic_decoderInterrupt_buffer_targetPrivilege;
  reg        [1:0]    PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped;
  reg        [3:0]    PrivilegedPlugin_logic_exception_code;
  wire                when_PrivilegedPlugin_l689;
  wire                when_PrivilegedPlugin_l702;
  wire                when_PrivilegedPlugin_l702_1;
  wire                when_PrivilegedPlugin_l702_2;
  wire                when_PrivilegedPlugin_l702_3;
  wire                when_PrivilegedPlugin_l702_4;
  wire                when_PrivilegedPlugin_l702_5;
  wire                when_PrivilegedPlugin_l702_6;
  wire       [1:0]    PrivilegedPlugin_logic_exception_targetPrivilege;
  wire                PrivilegedPlugin_logic_fsm_wantExit;
  reg                 PrivilegedPlugin_logic_fsm_wantStart;
  wire                PrivilegedPlugin_logic_fsm_wantKill;
  reg                 PrivilegedPlugin_logic_fsm_trap_fire;
  reg                 PrivilegedPlugin_logic_fsm_trap_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_fsm_trap_code;
  reg        [1:0]    PrivilegedPlugin_logic_fsm_trap_targetPrivilege;
  wire       [1:0]    PrivilegedPlugin_logic_fsm_xret_sourcePrivilege;
  reg        [1:0]    PrivilegedPlugin_logic_fsm_xret_targetPrivilege;
  wire                FetchPlugin_stages_0_haltRequest_PrivilegedPlugin_l968;
  wire                trap_fire /* verilator public */ ;
  wire       [3:0]    trap_code /* verilator public */ ;
  wire                trap_interrupt /* verilator public */ ;
  wire       [31:0]   trap_tval /* verilator public */ ;
  reg                 PerformanceCounterPlugin_logic_fsm_done;
  reg        [63:0]   PerformanceCounterPlugin_logic_fsm_resultCsr;
  reg        [63:0]   PerformanceCounterPlugin_logic_fsm_result;
  reg        [63:0]   PerformanceCounterPlugin_logic_fsm_ramReaded;
  reg        [5:0]    PerformanceCounterPlugin_logic_fsm_counterReaded;
  wire       [63:0]   PerformanceCounterPlugin_logic_fsm_calc;
  wire       [6:0]    PerformanceCounterPlugin_logic_flusher_hits;
  wire                PerformanceCounterPlugin_logic_flusher_hit;
  wire       [6:0]    PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input;
  wire       [6:0]    PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked;
  wire       [6:0]    PerformanceCounterPlugin_logic_flusher_oh;
  wire                _zz_PerformanceCounterPlugin_logic_flusher_sel;
  wire                _zz_PerformanceCounterPlugin_logic_flusher_sel_1;
  wire                _zz_PerformanceCounterPlugin_logic_flusher_sel_2;
  wire                _zz_PerformanceCounterPlugin_logic_flusher_sel_3;
  wire                _zz_PerformanceCounterPlugin_logic_flusher_sel_4;
  wire                _zz_PerformanceCounterPlugin_logic_flusher_sel_5;
  wire       [2:0]    PerformanceCounterPlugin_logic_flusher_sel;
  reg                 PerformanceCounterPlugin_logic_csrRead_fired;
  wire                PerformanceCounterPlugin_logic_fsm_csrReadCmd_fire;
  reg                 PerformanceCounterPlugin_logic_csrRead_requested;
  wire                when_PerformanceCounterPlugin_l253;
  reg                 PerformanceCounterPlugin_logic_csrWrite_fired;
  wire                PerformanceCounterPlugin_logic_fsm_csrWriteCmd_fire;
  wire                when_PerformanceCounterPlugin_l268;
  wire                when_MmuPlugin_l326;
  reg                 FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg;
  wire                when_MmuPlugin_l260_2;
  wire       [4:0]    FetchCachePlugin_logic_translationPort_logic_read_0_readAddress;
  wire       [41:0]   _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid;
  wire       [41:0]   _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid;
  wire       [41:0]   _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid;
  wire       [41:0]   _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid;
  wire       [4:0]    FetchCachePlugin_logic_translationPort_logic_read_1_readAddress;
  wire       [21:0]   _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid;
  wire       [21:0]   _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid;
  wire       [5:0]    FetchCachePlugin_logic_translationPort_logic_ctrl_hits;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hit;
  wire       [5:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_3;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_4;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_5;
  reg        [5:0]    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_1;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_2;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_3;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_4;
  wire       [5:0]    FetchCachePlugin_logic_translationPort_logic_ctrl_oh;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4;
  wire                _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineException;
  wire       [31:0]   FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault;
  reg                 FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_needRefill;
  wire                FetchCachePlugin_logic_translationPort_logic_ctrl_askRefill;
  wire                when_MmuPlugin_l297_1;
  wire                when_MmuPlugin_l298_1;
  wire                when_MmuPlugin_l326_1;
  wire                MmuPlugin_logic_refill_wantExit;
  reg                 MmuPlugin_logic_refill_wantStart;
  wire                MmuPlugin_logic_refill_wantKill;
  wire                MmuPlugin_logic_refill_busy;
  reg        [1:0]    MmuPlugin_logic_refill_portOhReg;
  wire                _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask;
  wire                _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask;
  reg        [31:0]   MmuPlugin_logic_refill_virtual;
  wire       [1:0]    MmuPlugin_logic_refill_portsRequests;
  reg                 MmuPlugin_logic_refill_portsRequest;
  wire       [1:0]    MmuPlugin_logic_refill_portsRequests_ohFirst_input;
  wire       [1:0]    MmuPlugin_logic_refill_portsRequests_ohFirst_masked;
  wire       [1:0]    MmuPlugin_logic_refill_portsOh;
  reg        [1:0]    MmuPlugin_logic_refill_portsOh_regNext;
  reg        [31:0]   _zz_MmuPlugin_logic_refill_portsAddress;
  reg        [31:0]   _zz_MmuPlugin_logic_refill_portsAddress_1;
  wire       [31:0]   MmuPlugin_logic_refill_portsAddress;
  reg        [1:0]    MmuPlugin_logic_refill_cacheRefill;
  reg                 MmuPlugin_logic_refill_cacheRefillAny;
  reg        [1:0]    MmuPlugin_logic_refill_cacheRefillSet;
  reg                 MmuPlugin_logic_refill_cacheRefillAnySet;
  wire                MmuPlugin_logic_refill_doWake;
  reg        [31:0]   MmuPlugin_logic_refill_load_address;
  reg                 MmuPlugin_logic_refill_load_rsp_valid;
  reg        [31:0]   MmuPlugin_logic_refill_load_rsp_payload_data;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_fault;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_redo;
  reg        [1:0]    MmuPlugin_logic_refill_load_rsp_payload_refillSlot;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_refillSlotAny;
  wire       [31:0]   MmuPlugin_logic_refill_load_readed;
  wire                when_MmuPlugin_l388;
  wire                MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_flags_R;
  wire                MmuPlugin_logic_refill_load_flags_W;
  wire                MmuPlugin_logic_refill_load_flags_X;
  wire                MmuPlugin_logic_refill_load_flags_U;
  wire                MmuPlugin_logic_refill_load_flags_G;
  wire                MmuPlugin_logic_refill_load_flags_A;
  wire                MmuPlugin_logic_refill_load_flags_D;
  wire       [31:0]   _zz_MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_leaf;
  reg                 MmuPlugin_logic_refill_load_exception;
  reg        [31:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_0;
  reg        [31:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_1;
  wire                MmuPlugin_logic_refill_load_levelException_0;
  reg                 MmuPlugin_logic_refill_load_levelException_1;
  reg        [31:0]   MmuPlugin_logic_refill_load_nextLevelBase;
  wire                when_MmuPlugin_l416;
  reg                 MmuPlugin_logic_invalidate_requested;
  reg                 MmuPlugin_logic_invalidate_canStart;
  reg        [5:0]    MmuPlugin_logic_invalidate_counter;
  wire                MmuPlugin_logic_invalidate_done;
  wire                when_MmuPlugin_l492;
  wire                FetchPlugin_stages_0_haltRequest_MmuPlugin_l503;
  wire                when_MmuPlugin_l505;
  wire                when_MmuPlugin_l511;
  reg                 MmuPlugin_logic_invalidate_done_regNext;
  wire                when_MmuPlugin_l515;
  wire                EU0_CsrAccessPlugin_logic_fsm_wantExit;
  reg                 EU0_CsrAccessPlugin_logic_fsm_wantStart;
  wire                EU0_CsrAccessPlugin_logic_fsm_wantKill;
  reg                 REG_CSR_773;
  reg                 REG_CSR_835;
  reg                 REG_CSR_833;
  reg                 REG_CSR_832;
  reg                 REG_CSR_3857;
  reg                 REG_CSR_3858;
  reg                 REG_CSR_3859;
  reg                 REG_CSR_3860;
  reg                 REG_CSR_769;
  reg                 REG_CSR_834;
  reg                 REG_CSR_768;
  reg                 REG_CSR_836;
  reg                 REG_CSR_772;
  reg                 REG_CSR_770;
  reg                 REG_CSR_771;
  reg                 REG_CSR_261;
  reg                 REG_CSR_323;
  reg                 REG_CSR_321;
  reg                 REG_CSR_320;
  reg                 REG_CSR_322;
  reg                 REG_CSR_256;
  reg                 REG_CSR_260;
  reg                 REG_CSR_324;
  reg                 REG_CSR_262;
  reg                 REG_CSR_774;
  reg                 REG_CSR_;
  reg                 REG_CSR_803;
  reg                 REG_CSR_804;
  reg                 REG_CSR_805;
  reg                 REG_CSR_806;
  reg                 REG_CSR_384;
  reg                 REG_CSR_PerformanceCounterPlugin_logic_csrFilter;
  wire                when_Pipeline_l278;
  reg                 Lsu2Plugin_logic_lqSqArbitration_s0_ready_output;
  wire                when_Pipeline_l278_1;
  wire                when_Connection_l74;
  reg        [8:0]    Lsu2Plugin_logic_special_atomic_stateReg;
  reg        [8:0]    Lsu2Plugin_logic_special_atomic_stateNext;
  wire                when_Lsu2Plugin_l1704;
  wire                when_Lsu2Plugin_l1705;
  wire                Lsu2Plugin_setup_cacheLoad_cmd_fire;
  wire                when_Lsu2Plugin_l1715;
  wire                when_Lsu2Plugin_l1824;
  wire                when_StateMachine_l253;
  wire                when_StateMachine_l253_1;
  reg        [2:0]    MmuPlugin_logic_refill_stateReg;
  reg        [2:0]    MmuPlugin_logic_refill_stateNext;
  wire                when_MmuPlugin_l452;
  wire                when_MmuPlugin_l452_1;
  wire                when_MmuPlugin_l461;
  wire                when_MmuPlugin_l469;
  wire                EU0_CsrAccessPlugin_logic_ramReadPort_valid;
  wire                EU0_CsrAccessPlugin_logic_ramReadPort_ready;
  wire       [4:0]    EU0_CsrAccessPlugin_logic_ramReadPort_address;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_ramReadPort_data;
  wire                EU0_CsrAccessPlugin_logic_ramWritePort_valid;
  wire                EU0_CsrAccessPlugin_logic_ramWritePort_ready;
  wire       [4:0]    EU0_CsrAccessPlugin_logic_ramWritePort_address;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_ramWritePort_data;
  reg        [5:0]    CsrRamPlugin_logic_flush_counter;
  wire                CsrRamPlugin_logic_flush_done;
  wire                when_CsrRamPlugin_l61;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_hits;
  wire                CsrRamPlugin_logic_writeLogic_hit;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_input;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_oh;
  wire                _zz_PerformanceCounterPlugin_setup_writePort_ready;
  wire                _zz_PrivilegedPlugin_setup_ramWrite_ready;
  wire                _zz_CsrRamPlugin_setup_initPort_ready;
  wire                _zz_CsrRamPlugin_logic_writeLogic_sel;
  wire                _zz_CsrRamPlugin_logic_writeLogic_sel_1;
  wire       [1:0]    CsrRamPlugin_logic_writeLogic_sel;
  wire                CsrRamPlugin_logic_writeLogic_port_valid;
  wire       [4:0]    CsrRamPlugin_logic_writeLogic_port_payload_address;
  wire       [31:0]   CsrRamPlugin_logic_writeLogic_port_payload_data;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_hits;
  wire                CsrRamPlugin_logic_readLogic_hit;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_input;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_oh;
  wire                _zz_PerformanceCounterPlugin_setup_readPort_ready;
  wire                _zz_PrivilegedPlugin_setup_ramRead_ready;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_sel;
  wire       [4:0]    CsrRamPlugin_logic_readLogic_port_address;
  wire       [31:0]   CsrRamPlugin_logic_readLogic_port_data;
  reg        [4:0]    EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_ramSel;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_regs_microOp;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_doImm;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_doMask;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_doClear;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_regs_rs1;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_implemented;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_trap;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_flushPipeline;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_read;
  reg                 EU0_CsrAccessPlugin_logic_fsm_regs_write;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_regs_aluInput;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_regs_csrValue;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_immZero;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_srcZero;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_csrWrite;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_csrRead;
  wire                COMB_CSR_773;
  wire                COMB_CSR_835;
  wire                COMB_CSR_833;
  wire                COMB_CSR_832;
  wire                COMB_CSR_3857;
  wire                COMB_CSR_3858;
  wire                COMB_CSR_3859;
  wire                COMB_CSR_3860;
  wire                COMB_CSR_769;
  wire                COMB_CSR_834;
  wire                COMB_CSR_768;
  wire                COMB_CSR_836;
  wire                COMB_CSR_772;
  wire                COMB_CSR_770;
  wire                COMB_CSR_771;
  wire                COMB_CSR_261;
  wire                COMB_CSR_323;
  wire                COMB_CSR_321;
  wire                COMB_CSR_320;
  wire                COMB_CSR_322;
  wire                COMB_CSR_256;
  wire                COMB_CSR_260;
  wire                COMB_CSR_324;
  wire                COMB_CSR_262;
  wire                COMB_CSR_774;
  wire                COMB_CSR_;
  wire                COMB_CSR_803;
  wire                COMB_CSR_804;
  wire                COMB_CSR_805;
  wire                COMB_CSR_806;
  wire                COMB_CSR_384;
  wire                COMB_CSR_PerformanceCounterPlugin_logic_csrFilter;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_trap;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_write;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_read;
  wire                EU0_CsrAccessPlugin_logic_fsm_startLogic_onDecodeDo;
  wire                when_CsrAccessPlugin_l181;
  reg                 EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  reg                 EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15;
  reg        [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16;
  wire                when_CsrAccessPlugin_l244;
  wire       [31:0]   _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17;
  reg        [31:0]   EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire                when_CsrAccessPlugin_l270;
  wire                when_CsrAccessPlugin_l276;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_masked;
  wire       [31:0]   EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
  reg                 EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  reg                 EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo;
  wire                when_CsrAccessPlugin_l326;
  wire                when_CsrAccessPlugin_l326_1;
  wire                when_CsrAccessPlugin_l326_2;
  wire                when_CsrAccessPlugin_l326_3;
  wire                when_CsrAccessPlugin_l326_4;
  wire                when_CsrAccessPlugin_l326_5;
  wire                when_CsrAccessPlugin_l326_6;
  wire                when_CsrAccessPlugin_l326_7;
  wire                when_CsrAccessPlugin_l326_8;
  wire                when_CsrAccessPlugin_l326_9;
  wire                when_CsrAccessPlugin_l326_10;
  wire                when_CsrAccessPlugin_l326_11;
  wire                when_CsrAccessPlugin_l326_12;
  wire                when_CsrAccessPlugin_l326_13;
  wire                when_CsrAccessPlugin_l331;
  wire                when_CsrAccessPlugin_l326_14;
  wire                when_CsrAccessPlugin_l325;
  wire                when_PerformanceCounterPlugin_l273;
  wire                when_PerformanceCounterPlugin_l275;
  reg                 EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired;
  wire                when_CsrAccessPlugin_l336;
  wire                when_CsrAccessPlugin_l340;
  reg                 EU0_CsrAccessPlugin_logic_fsm_isDone;
  reg                 EU0_CsrAccessPlugin_logic_fsm_isCompletionReady;
  reg        [2:0]    EU0_CsrAccessPlugin_logic_fsm_stateReg;
  reg        [2:0]    EU0_CsrAccessPlugin_logic_fsm_stateNext;
  wire       [11:0]   switch_CsrAccessPlugin_l204;
  wire                when_CsrAccessPlugin_l283;
  wire                when_CsrAccessPlugin_l309;
  wire                EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_CsrAccessPlugin_l373;
  wire                when_CsrAccessPlugin_l376;
  wire                csrAccess_valid /* verilator public */ ;
  wire       [5:0]    csrAccess_payload_robId /* verilator public */ ;
  wire       [11:0]   csrAccess_payload_address /* verilator public */ ;
  wire       [31:0]   csrAccess_payload_write /* verilator public */ ;
  wire       [31:0]   csrAccess_payload_read /* verilator public */ ;
  wire                csrAccess_payload_writeDone /* verilator public */ ;
  wire                csrAccess_payload_readDone /* verilator public */ ;
  wire                EU0_ExecutionUnitBase_pipeline_execute_2_isFireing;
  wire                DecoderPlugin_logic_slots_0_rdZero;
  wire                _zz_FrontendPlugin_decoded_SQ_ALLOC_0;
  wire                _zz_FrontendPlugin_decoded_SQ_ALLOC_0_1;
  reg                 DecoderPlugin_logic_slots_0_x0AlwaysZero;
  wire                _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_0;
  wire                _zz_FrontendPlugin_decoded_WRITE_RD_0;
  wire                _zz_FrontendPlugin_decoded_IS_ANY_0;
  wire                DecoderPlugin_logic_slots_1_rdZero;
  wire                _zz_FrontendPlugin_decoded_SQ_ALLOC_1;
  wire                _zz_FrontendPlugin_decoded_SQ_ALLOC_1_1;
  reg                 DecoderPlugin_logic_slots_1_x0AlwaysZero;
  wire                _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_1;
  wire                _zz_FrontendPlugin_decoded_IS_JAL_1;
  wire                _zz_FrontendPlugin_decoded_IS_ANY_1;
  wire                DecoderPlugin_logic_exception_set;
  wire                DecoderPlugin_logic_exception_clear;
  reg                 DecoderPlugin_logic_exception_trigged;
  wire                when_DecoderPlugin_l302;
  reg                 DecoderPlugin_logic_exception_exceptionReg_0;
  reg                 DecoderPlugin_logic_exception_exceptionReg_1;
  wire                when_DecoderPlugin_l303;
  reg                 DecoderPlugin_logic_exception_fetchFaultReg_0;
  reg                 DecoderPlugin_logic_exception_fetchFaultReg_1;
  wire                when_DecoderPlugin_l304;
  reg                 DecoderPlugin_logic_exception_fetchFaultPageReg_0;
  reg                 DecoderPlugin_logic_exception_fetchFaultPageReg_1;
  wire                when_DecoderPlugin_l306;
  reg                 DecoderPlugin_logic_exception_debugEnterReg_0;
  reg                 DecoderPlugin_logic_exception_debugEnterReg_1;
  wire                when_DecoderPlugin_l307;
  reg        [31:0]   DecoderPlugin_logic_exception_epcReg_0;
  reg        [31:0]   DecoderPlugin_logic_exception_epcReg_1;
  wire                when_DecoderPlugin_l308;
  reg        [31:0]   DecoderPlugin_logic_exception_instReg_0;
  reg        [31:0]   DecoderPlugin_logic_exception_instReg_1;
  wire       [1:0]    _zz_DecoderPlugin_setup_exceptionPort_payload_tval;
  wire                _zz_DecoderPlugin_setup_exceptionPort_payload_tval_1;
  wire                DecoderPlugin_logic_exception_fetchFault;
  wire                DecoderPlugin_logic_exception_fetchFaultPage;
  wire                DecoderPlugin_logic_exception_debugEnter;
  wire       [31:0]   DecoderPlugin_logic_exception_pc;
  wire                DecoderPlugin_logic_exception_pipelineEmpty;
  wire                DecoderPlugin_logic_exception_doIt;
  reg                 DecoderPlugin_logic_exception_doItAgain;
  wire                _zz_FrontendPlugin_decoded_isFlushingRoot;
  wire                FrontendPlugin_decoded_haltRequest_DecoderPlugin_l322;
  wire                FrontendPlugin_decoded_haltRequest_DecoderPlugin_l323;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_1;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_1;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_1;
  wire                _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_1;
  wire                switch_Misc_l232_3;
  reg        [31:0]   _zz_FrontendPlugin_decoded_OFFSET_0;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rs1Link;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdEquRs1;
  wire       [1:0]    DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_0_applyIt_badTaken;
  wire                when_DecoderPredictionPlugin_l212;
  wire                when_DecoderPredictionPlugin_l213;
  wire                when_DecoderPredictionPlugin_l219;
  wire                switch_Misc_l232_4;
  reg        [31:0]   _zz_FrontendPlugin_decoded_OFFSET_1;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rdLink;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rs1Link;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rdEquRs1;
  wire       [1:0]    DecoderPredictionPlugin_logic_decodePatch_slots_1_pcAdd_slices;
  wire                DecoderPredictionPlugin_logic_decodePatch_slots_1_applyIt_badTaken;
  wire                when_DecoderPredictionPlugin_l212_1;
  wire                when_DecoderPredictionPlugin_l213_1;
  wire                when_DecoderPredictionPlugin_l219_1;
  wire                DecoderPredictionPlugin_logic_decodePatch_applyIt_hit;
  wire                FrontendPlugin_serialized_isFireing;
  reg                 DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle;
  wire                when_DecoderPredictionPlugin_l236;
  wire                when_DecoderPredictionPlugin_l243;
  wire                when_DecoderPredictionPlugin_l244;
  wire                ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address;
  reg        [31:0]   ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                ALU0_ExecutionUnitBase_pipeline_push_port_valid;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_push_port_robId;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_push_port_physRd;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1;
  wire       [1:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2;
  wire                ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  wire       [31:0]   ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId;
  wire                ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  wire                ALU0_ExecutionUnitBase_pipeline_execute_0_isFireing;
  wire                ALU0_ExecutionUnitBase_pipeline_completion_1_port_valid;
  wire       [5:0]    ALU0_ExecutionUnitBase_pipeline_completion_1_port_payload_id;
  wire                ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address;
  reg        [31:0]   ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                ALU1_ExecutionUnitBase_pipeline_push_port_valid;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_push_port_robId;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_push_port_physRd;
  wire                _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2;
  wire                _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1;
  wire       [1:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2;
  wire                ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_valid;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  wire       [31:0]   ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_robId;
  wire                ALU1_ExecutionUnitBase_pipeline_completion_0_port_valid;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  wire                ALU1_ExecutionUnitBase_pipeline_execute_0_isFireing;
  wire                ALU1_ExecutionUnitBase_pipeline_completion_1_port_valid;
  wire       [5:0]    ALU1_ExecutionUnitBase_pipeline_completion_1_port_payload_id;
  wire                EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address;
  reg        [31:0]   EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                EU0_ExecutionUnitBase_pipeline_push_port_valid;
  wire                EU0_ExecutionUnitBase_pipeline_push_port_ready;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_push_port_robId;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_push_port_physRd;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_push_port_context_0;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_push_port_context_1;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD;
  wire                EU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid;
  wire                EU0_ExecutionUnitBase_pipeline_writeBack_0_write_ready;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  wire       [31:0]   EU0_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId;
  wire                EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_ExecutionUnitBase_l303;
  wire                EU0_ExecutionUnitBase_pipeline_completion_0_port_valid;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  wire                EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_fire;
  wire                EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_valid;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_payload_robId;
  wire                EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_fire;
  wire                EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_valid;
  wire       [5:0]    EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_payload_physical;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_1_ready_output;
  reg                 EU0_ExecutionUnitBase_pipeline_execute_0_ready_output;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_1_ready_output;
  wire                EU0_ExecutionUnitBase_pipeline_fetch_1_ready;
  reg                 EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output;
  wire                when_Pipeline_l278_2;
  wire                when_Pipeline_l278_3;
  wire                when_Pipeline_l278_4;
  wire                when_Connection_l74_1;
  wire                when_Connection_l74_2;
  wire                when_Connection_l74_3;
  wire                BranchContextPlugin_free_dispatchMem_writes_0_port_valid;
  wire       [3:0]    BranchContextPlugin_free_dispatchMem_writes_0_port_payload_address;
  wire       [28:0]   BranchContextPlugin_free_dispatchMem_writes_0_port_payload_data;
  wire                BranchContextPlugin_free_dispatchMem_writes_1_port_valid;
  wire       [3:0]    BranchContextPlugin_free_dispatchMem_writes_1_port_payload_address;
  wire       [28:0]   BranchContextPlugin_free_dispatchMem_writes_1_port_payload_data;
  wire                BranchContextPlugin_free_learn_valid;
  wire       [3:0]    BranchContextPlugin_free_learn_bid;
  wire       [64:0]   _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice;
  wire       [28:0]   BranchContextPlugin_free_learn_raw;
  wire       [3:0]    _zz_BranchContextPlugin_free_learn_GSHARE_COUNTER_0;
  wire       [31:0]   DispatchPlugin_logic_queueStaticWakeTransposed_0;
  wire       [31:0]   DispatchPlugin_logic_queueStaticWakeTransposedHistory_0_0;
  reg        [5:0]    DispatchPlugin_logic_ptr_next;
  reg        [5:0]    DispatchPlugin_logic_ptr_current;
  wire                toplevel_DispatchPlugin_logic_queue_io_push_fire;
  wire                FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l187;
  wire                DispatchPlugin_logic_push_skip;
  wire                DispatchPlugin_logic_push_fenceOlder;
  wire                DispatchPlugin_logic_push_fenceYounger;
  wire                when_DispatchPlugin_l192;
  reg                 DispatchPlugin_logic_push_fenceYoungerLast;
  wire                DispatchPlugin_logic_push_commitNotWaitingOnUs;
  wire                FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l195;
  wire                FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l196;
  wire       [31:0]   DispatchPlugin_logic_push_slots_0_self;
  wire       [31:0]   DispatchPlugin_logic_push_slots_0_events_0;
  wire       [31:0]   DispatchPlugin_logic_push_slots_0_events_1;
  wire       [31:0]   DispatchPlugin_logic_push_slots_1_self;
  wire       [31:0]   DispatchPlugin_logic_push_slots_1_events_0;
  wire       [31:0]   DispatchPlugin_logic_push_slots_1_events_1;
  wire                DispatchPlugin_logic_pop_0_stagesList_0_valid;
  reg                 DispatchPlugin_logic_pop_0_stagesList_1_valid;
  wire       [31:0]   DispatchPlugin_logic_pop_0_portEventFull;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_1;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_2;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_4;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_5;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_6;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_7;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_8;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_9;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_10;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_11;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_12;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_13;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_14;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_15;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_16;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_17;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_18;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_19;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_20;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_21;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_22;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_23;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_24;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_25;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_26;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_27;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_28;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_29;
  wire                _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_30;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_4;
  wire                toplevel_DispatchPlugin_logic_queue_io_schedules_0_fire;
  wire       [31:0]   DispatchPlugin_logic_pop_0_wake_L0_mask;
  wire                DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid;
  wire       [5:0]    DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical;
  wire                DispatchPlugin_logic_pop_1_stagesList_0_valid;
  reg                 DispatchPlugin_logic_pop_1_stagesList_1_valid;
  wire       [31:0]   DispatchPlugin_logic_pop_1_portEventFull;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_1;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_2;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_4;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_5;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_6;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_7;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_8;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_9;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_10;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_11;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_12;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_13;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_14;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_15;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_16;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_17;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_18;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_19;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_20;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_21;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_22;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_23;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_24;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_25;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_26;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_27;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_28;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_29;
  wire                _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_30;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_0;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_1;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_2;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_3;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_4;
  wire                toplevel_DispatchPlugin_logic_queue_io_schedules_1_fire;
  wire       [31:0]   DispatchPlugin_logic_pop_1_wake_L0_mask;
  wire                DispatchPlugin_logic_pop_1_wake_L0_bypassed_valid;
  wire       [5:0]    DispatchPlugin_logic_pop_1_wake_L0_bypassed_payload_physical;
  wire                DispatchPlugin_logic_pop_2_stagesList_0_valid;
  reg                 DispatchPlugin_logic_pop_2_stagesList_1_valid;
  wire       [31:0]   DispatchPlugin_logic_pop_2_portEventFull;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_1;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_2;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_3;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_4;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_5;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_6;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_7;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_8;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_9;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_10;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_11;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_12;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_13;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_14;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_15;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_16;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_17;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_18;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_19;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_20;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_21;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_22;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_23;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_24;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_25;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_26;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_27;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_28;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_29;
  wire                _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_30;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_0;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_1;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_2;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_3;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_4;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_5;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_6;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_7;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_8;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_9;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_10;
  wire                DispatchPlugin_logic_pop_2_stagesList_1_haltRequest_DispatchPlugin_l292;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_0;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_1;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_2;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_3;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_4;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_5;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_6;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_7;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_8;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_9;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_10;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_0;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_1;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_2;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_3;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_4;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_5;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_6;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_7;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_8;
  wire       [2:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_9;
  wire       [1:0]    _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_10;
  reg                 DispatchPlugin_logic_pop_2_stagesList_0_ready_output;
  wire                when_Pipeline_l278_5;
  wire                when_Connection_l74_4;
  wire                DispatchPlugin_logic_wake_dynamic_offseted_0_valid;
  wire       [4:0]    DispatchPlugin_logic_wake_dynamic_offseted_0_payload;
  wire                DispatchPlugin_logic_wake_dynamic_offseted_1_valid;
  wire       [4:0]    DispatchPlugin_logic_wake_dynamic_offseted_1_payload;
  wire                DispatchPlugin_logic_wake_dynamic_offseted_2_valid;
  wire       [4:0]    DispatchPlugin_logic_wake_dynamic_offseted_2_payload;
  wire                DispatchPlugin_logic_wake_dynamic_offseted_3_valid;
  wire       [4:0]    DispatchPlugin_logic_wake_dynamic_offseted_3_payload;
  wire       [31:0]   DispatchPlugin_logic_wake_dynamic_masks_0;
  wire       [31:0]   DispatchPlugin_logic_wake_dynamic_masks_1;
  wire       [31:0]   DispatchPlugin_logic_wake_dynamic_masks_2;
  wire       [31:0]   DispatchPlugin_logic_wake_dynamic_masks_3;
  wire       [31:0]   DispatchPlugin_logic_wake_statics_0_popMask;
  wire       [31:0]   DispatchPlugin_logic_wake_statics_0_history_0;
  (* keep , syn_keep *) wire       [31:0]   DispatchPlugin_logic_wake_optReduce_relaxed /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   DispatchPlugin_logic_wake_optReduce_reduced;
  wire                DispatchPlugin_logic_whitebox_issuePorts_0_valid /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_0_payload_robId /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_0_payload_physRd /* verilator public */ ;
  wire                DispatchPlugin_logic_whitebox_issuePorts_1_valid /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_1_payload_robId /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_1_payload_physRd /* verilator public */ ;
  wire                DispatchPlugin_logic_whitebox_issuePorts_2_valid /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_2_payload_robId /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_2_payload_physRd /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_2_payload_context_0 /* verilator public */ ;
  wire       [5:0]    DispatchPlugin_logic_whitebox_issuePorts_2_payload_context_1 /* verilator public */ ;
  wire                integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_0_bus_robId;
  wire                integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data;
  wire                integer_RegFilePlugin_logic_writeMerges_1_bus_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_1_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_1_bus_data;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_1_bus_robId;
  wire                integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data;
  wire                integer_RegFilePlugin_logic_writeMerges_2_bus_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_2_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_2_bus_data;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_2_bus_robId;
  wire                integer_RegFilePlugin_logic_writeMerges_2_bypass_port_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_2_bypass_port_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_2_bypass_port_data;
  wire                integer_RegFilePlugin_logic_writeMerges_3_bus_valid;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_3_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_3_bus_data;
  wire       [5:0]    integer_RegFilePlugin_logic_writeMerges_3_bus_robId;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1;
  wire                when_RegFilePlugin_l322;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1;
  wire                when_RegFilePlugin_l322_1;
  wire                _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1;
  wire                when_RegFilePlugin_l322_2;
  wire                _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1;
  wire                when_RegFilePlugin_l322_3;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1;
  wire                when_RegFilePlugin_l322_4;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  wire                _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1;
  wire                when_RegFilePlugin_l322_5;
  wire                integer_write_0_valid /* verilator public */ ;
  wire       [5:0]    integer_write_0_address /* verilator public */ ;
  wire       [31:0]   integer_write_0_data /* verilator public */ ;
  wire       [5:0]    integer_write_0_robId /* verilator public */ ;
  wire                integer_write_1_valid /* verilator public */ ;
  wire       [5:0]    integer_write_1_address /* verilator public */ ;
  wire       [31:0]   integer_write_1_data /* verilator public */ ;
  wire       [5:0]    integer_write_1_robId /* verilator public */ ;
  wire                integer_write_2_valid /* verilator public */ ;
  wire       [5:0]    integer_write_2_address /* verilator public */ ;
  wire       [31:0]   integer_write_2_data /* verilator public */ ;
  wire       [5:0]    integer_write_2_robId /* verilator public */ ;
  wire                integer_write_3_valid /* verilator public */ ;
  wire       [5:0]    integer_write_3_address /* verilator public */ ;
  wire       [31:0]   integer_write_3_data /* verilator public */ ;
  wire       [5:0]    integer_write_3_robId /* verilator public */ ;
  wire                RobPlugin_logic_completionMem_targetWrite_valid;
  wire       [4:0]    RobPlugin_logic_completionMem_targetWrite_payload_address;
  reg        [1:0]    RobPlugin_logic_completionMem_targetWrite_payload_data;
  wire       [5:0]    RobPlugin_logic_completionMem_init_0_robId;
  wire       [5:0]    RobPlugin_logic_completionMem_init_1_robId;
  wire       [4:0]    RobPlugin_logic_completionMem_reads_0_targetRead_address;
  wire       [1:0]    RobPlugin_logic_completionMem_reads_0_targetRead_data;
  wire       [5:0]    _zz_CommitPlugin_setup_robLineMask_mask;
  wire       [5:0]    _zz_CommitPlugin_setup_robLineMask_mask_1;
  wire       [5:0]    _zz_when_RobPlugin_l118;
  wire                when_RobPlugin_l118;
  wire                when_RobPlugin_l118_1;
  wire                when_RobPlugin_l118_2;
  wire                when_RobPlugin_l118_3;
  wire                when_RobPlugin_l118_4;
  wire                when_RobPlugin_l118_5;
  wire                when_RobPlugin_l118_6;
  wire       [5:0]    _zz_when_RobPlugin_l118_1;
  wire                when_RobPlugin_l118_7;
  wire                when_RobPlugin_l118_8;
  wire                when_RobPlugin_l118_9;
  wire                when_RobPlugin_l118_10;
  wire                when_RobPlugin_l118_11;
  wire                when_RobPlugin_l118_12;
  wire                when_RobPlugin_l118_13;
  wire                when_RobPlugin_l123;
  wire       [4:0]    _zz_CommitPlugin_logic_commit_active;
  wire       [1:0]    _zz_CommitPlugin_logic_commit_active_1;
  wire       [1:0]    _zz_CommitPlugin_logic_commit_active_2;
  wire       [4:0]    _zz_integer_RfAllocationPlugin_logic_push_mask_0;
  wire       [1:0]    _zz_integer_RfAllocationPlugin_logic_push_mask_0_1;
  wire       [1:0]    _zz_integer_RfAllocationPlugin_logic_push_mask_0_2;
  wire       [4:0]    _zz_224;
  wire       [4:0]    _zz_commit_pc_0;
  wire       [63:0]   _zz_commit_pc_0_1;
  wire       [4:0]    _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc;
  wire       [63:0]   _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_1;
  wire       [4:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire       [4:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  wire       [63:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_1;
  wire       [4:0]    _zz_235;
  wire       [4:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0;
  wire       [1:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1;
  wire       [4:0]    _zz_integer_RfAllocationPlugin_logic_push_writeRd_0;
  wire       [1:0]    _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1;
  wire       [4:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire       [4:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1;
  wire       [4:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0;
  wire       [11:0]   _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_1;
  wire       [11:0]   _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2;
  wire       [4:0]    _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0;
  wire       [11:0]   _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_1;
  wire       [11:0]   _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2;
  wire       [4:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0;
  wire       [9:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_1;
  wire       [9:0]    _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2;
  wire       [4:0]    _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0;
  wire       [11:0]   _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_1;
  wire       [11:0]   _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2;
  wire       [4:0]    _zz_BranchContextPlugin_logic_onCommit_isBranch_0;
  wire       [1:0]    _zz_BranchContextPlugin_logic_onCommit_isBranch_0_1;
  wire       [1:0]    _zz_BranchContextPlugin_logic_onCommit_isBranch_0_2;
  wire       [4:0]    _zz_255;
  wire       [4:0]    _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0;
  wire       [1:0]    _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1;
  wire       [4:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch;
  wire       [1:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_1;
  wire       [4:0]    _zz_io_read_0_cmd_payload;
  wire       [1:0]    _zz_HistoryPlugin_logic_onCommit_isTaken_0;
  wire       [4:0]    _zz_262;
  wire       [4:0]    _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory;
  wire       [47:0]   _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_1;
  wire       [4:0]    _zz_267;
  wire       [4:0]    _zz_DecoderPredictionPlugin_logic_ras_healPush;
  wire       [7:0]    _zz_DecoderPredictionPlugin_logic_ras_healPush_1;
  wire       [4:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0;
  wire       [1:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_1;
  wire       [1:0]    _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2;
  wire       [4:0]    _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_1;
  wire       [1:0]    _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2;
  wire       [4:0]    _zz_276;
  wire       [4:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  wire       [4:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
  wire       [63:0]   _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1;
  wire       [4:0]    _zz_283;
  wire       [4:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  wire       [4:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  wire       [4:0]    _zz_288;
  wire       [4:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [4:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1;
  wire       [4:0]    _zz_295;
  wire       [4:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  wire       [4:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  wire       [4:0]    _zz_300;
  wire       [4:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire       [4:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1;
  wire       [4:0]    _zz_307;
  wire       [4:0]    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID;
  wire       [4:0]    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID;
  wire       [4:0]    _zz_312;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID;
  wire       [9:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_1;
  wire       [4:0]    _zz_317;
  wire       [4:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB;
  wire       [1:0]    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_1;
  wire                RobPlugin_logic_whitebox_completionsPorts_0_valid /* verilator public */ ;
  wire       [5:0]    RobPlugin_logic_whitebox_completionsPorts_0_payload_id /* verilator public */ ;
  wire                RobPlugin_logic_whitebox_completionsPorts_1_valid /* verilator public */ ;
  wire       [5:0]    RobPlugin_logic_whitebox_completionsPorts_1_payload_id /* verilator public */ ;
  wire                RobPlugin_logic_whitebox_completionsPorts_2_valid /* verilator public */ ;
  wire       [5:0]    RobPlugin_logic_whitebox_completionsPorts_2_payload_id /* verilator public */ ;
  wire                RobPlugin_logic_whitebox_completionsPorts_3_valid /* verilator public */ ;
  wire       [5:0]    RobPlugin_logic_whitebox_completionsPorts_3_payload_id /* verilator public */ ;
  wire                RobPlugin_logic_whitebox_completionsPorts_4_valid /* verilator public */ ;
  wire       [5:0]    RobPlugin_logic_whitebox_completionsPorts_4_payload_id /* verilator public */ ;
  wire                RobPlugin_logic_whitebox_completionsPorts_5_valid /* verilator public */ ;
  wire       [5:0]    RobPlugin_logic_whitebox_completionsPorts_5_payload_id /* verilator public */ ;
  wire                RobPlugin_logic_whitebox_completionsPorts_6_valid /* verilator public */ ;
  wire       [5:0]    RobPlugin_logic_whitebox_completionsPorts_6_payload_id /* verilator public */ ;
  reg        [6:0]    RfDependencyPlugin_logic_forRf_integer_init_counter;
  wire                RfDependencyPlugin_logic_forRf_integer_init_busy;
  reg                 _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0;
  reg        [5:0]    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0;
  wire                when_RfDependencyPlugin_l241;
  wire                when_RfDependencyPlugin_l241_1;
  wire                when_RfDependencyPlugin_l245;
  reg                 _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0;
  reg        [5:0]    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0;
  wire                when_RfDependencyPlugin_l241_2;
  wire                when_RfDependencyPlugin_l241_3;
  wire                when_RfDependencyPlugin_l245_1;
  reg                 _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1;
  reg        [5:0]    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_1;
  wire                when_RfDependencyPlugin_l235;
  wire                when_RfDependencyPlugin_l241_4;
  wire                when_RfDependencyPlugin_l241_5;
  wire                when_RfDependencyPlugin_l245_2;
  reg                 _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1;
  reg        [5:0]    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_1;
  wire                when_RfDependencyPlugin_l235_1;
  wire                when_RfDependencyPlugin_l241_6;
  wire                when_RfDependencyPlugin_l241_7;
  wire                when_RfDependencyPlugin_l245_3;
  reg                 FrontendPlugin_allocated_ready_output;
  wire                FrontendPlugin_serialized_ready_output;
  wire                when_Connection_l66;
  reg                 FrontendPlugin_decoded_ready_output;
  wire                _zz_FrontendPlugin_decompressed_isFlushed;
  wire                FrontendPlugin_decompressed_ready_output;
  wire                FrontendPlugin_decompressed_ready;
  wire                FrontendPlugin_aligned_ready_output;
  wire                when_Pipeline_l278_6;
  wire                when_Pipeline_l285;
  wire                when_Pipeline_l278_7;
  wire                when_Pipeline_l278_8;
  wire                when_Connection_l74_5;
  wire                when_Connection_l74_6;
  reg        [6:0]    PcPlugin_logic_init_counter;
  wire                PcPlugin_logic_init_booted;
  wire                PcPlugin_logic_fetchPc_output_valid;
  wire                PcPlugin_logic_fetchPc_output_ready;
  wire       [31:0]   PcPlugin_logic_fetchPc_output_payload;
  reg        [31:0]   PcPlugin_logic_fetchPc_pcReg /* verilator public */ ;
  reg                 PcPlugin_logic_fetchPc_correction;
  reg                 PcPlugin_logic_fetchPc_correctionReg;
  wire                PcPlugin_logic_fetchPc_output_fire;
  wire                PcPlugin_logic_fetchPc_corrected;
  wire                PcPlugin_logic_fetchPc_pcRegPropagate;
  reg                 PcPlugin_logic_fetchPc_inc;
  wire                when_PcPlugin_l82;
  wire                when_PcPlugin_l82_1;
  reg        [31:0]   PcPlugin_logic_fetchPc_pc;
  reg                 PcPlugin_logic_fetchPc_flushed;
  wire                when_PcPlugin_l98;
  wire                PcPlugin_logic_fetchPc_fetcherHalt;
  wire                fetchLastFire /* verilator public */ ;
  wire       [11:0]   fetchLastId /* verilator public */ ;
  wire                FetchPlugin_stages_2_ready_output;
  wire                when_Connection_l66_1;
  reg                 FetchPlugin_stages_1_ready_output;
  wire                when_Connection_l54;
  reg                 FetchPlugin_stages_0_ready_output;
  wire                when_Pipeline_l278_9;
  wire                when_Pipeline_l278_10;
  wire                when_Connection_l74_7;
  wire                when_Connection_l74_8;
  reg                 FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid;
  reg        [63:0]   FetchPlugin_stages_2_Fetch_WORD_s2mBuffer;
  reg        [31:0]   FetchPlugin_stages_2_Fetch_FETCH_PC_s2mBuffer;
  reg                 FetchPlugin_stages_2_Fetch_WORD_FAULT_s2mBuffer;
  reg                 FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE_s2mBuffer;
  reg        [23:0]   FetchPlugin_stages_2_BRANCH_HISTORY_s2mBuffer;
  reg        [11:0]   FetchPlugin_stages_2_FETCH_ID_s2mBuffer;
  reg        [0:0]    FetchPlugin_stages_2_Prediction_WORD_BRANCH_SLICE_s2mBuffer;
  reg                 FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID_s2mBuffer;
  reg        [1:0]    FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT_s2mBuffer;
  reg        [31:0]   FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT_s2mBuffer;
  reg                 FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID_s2mBuffer;
  reg        [0:0]    FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_SLICE_s2mBuffer;
  reg                 FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE_s2mBuffer;
  reg        [1:0]    FetchPlugin_stages_2_GSHARE_COUNTER_s2mBuffer_0;
  reg        [1:0]    FetchPlugin_stages_2_GSHARE_COUNTER_s2mBuffer_1;
  reg        [31:0]   FetchPlugin_stages_2_Fetch_FETCH_PC_INC_s2mBuffer;
  reg        [3:0]    PerformanceCounterPlugin_logic_fsm_stateReg;
  reg        [3:0]    PerformanceCounterPlugin_logic_fsm_stateNext;
  wire                when_PerformanceCounterPlugin_l201;
  wire                when_PerformanceCounterPlugin_l161;
  wire                when_PerformanceCounterPlugin_l169;
  reg        [3:0]    PrivilegedPlugin_logic_fsm_stateReg;
  reg        [3:0]    PrivilegedPlugin_logic_fsm_stateNext;
  wire                when_PrivilegedPlugin_l766;
  reg        [4:0]    _zz_PrivilegedPlugin_setup_ramWrite_address;
  reg        [4:0]    _zz_PrivilegedPlugin_setup_ramWrite_address_1;
  reg        [4:0]    _zz_PrivilegedPlugin_setup_ramRead_address;
  reg        [4:0]    _zz_PrivilegedPlugin_setup_ramRead_address_1;
  wire                when_PrivilegedPlugin_l952;
  wire       [1:0]    switch_PrivilegedPlugin_l953;
  wire                when_StateMachine_l253_2;
  reg        [63:0]   _zz_FetchCachePlugin_logic_banks_0_read_rsp;
  reg                 when_MultiportRam_l328;
  reg        [63:0]   _zz_FetchCachePlugin_logic_banks_1_read_rsp;
  reg                 when_MultiportRam_l328_1;
  reg        [63:0]   _zz_FetchCachePlugin_logic_banks_2_read_rsp;
  reg                 when_MultiportRam_l328_2;
  reg        [63:0]   _zz_FetchCachePlugin_logic_banks_3_read_rsp;
  reg                 when_MultiportRam_l328_3;
  reg        [3:0]    _zz_FetchPlugin_stages_1_GSHARE_COUNTER_0_1;
  reg                 when_MultiportRam_l328_4;
  reg        [22:0]   _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_2;
  reg                 when_MultiportRam_l362;
  reg        [22:0]   _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_3;
  reg        [5:0]    _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter_1;
  reg                 when_MultiportRam_l362_1;
  reg        [5:0]    _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter_2;
  `ifndef SYNTHESIS
  reg [31:0] ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string;
  reg [63:0] ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string;
  reg [39:0] ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [31:0] ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string;
  reg [39:0] ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [63:0] ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string;
  reg [31:0] ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string;
  reg [63:0] ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string;
  reg [39:0] ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [31:0] ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string;
  reg [39:0] ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [63:0] ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string;
  reg [31:0] ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string;
  reg [31:0] ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string;
  reg [87:0] Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string;
  reg [87:0] Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string;
  reg [31:0] ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string;
  reg [63:0] ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string;
  reg [39:0] ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [31:0] ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string;
  reg [63:0] ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string;
  reg [39:0] ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [119:0] EnvCallPlugin_logic_flushes_stateReg_string;
  reg [119:0] EnvCallPlugin_logic_flushes_stateNext_string;
  reg [79:0] Lsu2Plugin_logic_special_atomic_stateReg_string;
  reg [79:0] Lsu2Plugin_logic_special_atomic_stateNext_string;
  reg [39:0] MmuPlugin_logic_refill_stateReg_string;
  reg [39:0] MmuPlugin_logic_refill_stateNext_string;
  reg [39:0] EU0_CsrAccessPlugin_logic_fsm_stateReg_string;
  reg [39:0] EU0_CsrAccessPlugin_logic_fsm_stateNext_string;
  reg [63:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string;
  reg [63:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string;
  reg [63:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string;
  reg [39:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string;
  reg [39:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string;
  reg [31:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string;
  reg [31:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string;
  reg [31:0] _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string;
  reg [63:0] _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string;
  reg [63:0] _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string;
  reg [63:0] _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string;
  reg [39:0] _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string;
  reg [39:0] _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string;
  reg [31:0] _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string;
  reg [31:0] _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string;
  reg [31:0] _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string;
  reg [159:0] PerformanceCounterPlugin_logic_fsm_stateReg_string;
  reg [159:0] PerformanceCounterPlugin_logic_fsm_stateNext_string;
  reg [79:0] PrivilegedPlugin_logic_fsm_stateReg_string;
  reg [79:0] PrivilegedPlugin_logic_fsm_stateNext_string;
  `endif

  reg [63:0] FetchCachePlugin_logic_banks_0_mem [0:511];
  reg [63:0] FetchCachePlugin_logic_banks_1_mem [0:511];
  reg [63:0] FetchCachePlugin_logic_banks_2_mem [0:511];
  reg [63:0] FetchCachePlugin_logic_banks_3_mem [0:511];
  (* ram_style = "distributed" *) reg [21:0] FetchCachePlugin_logic_ways_0_mem [0:63];
  (* ram_style = "distributed" *) reg [21:0] FetchCachePlugin_logic_ways_1_mem [0:63];
  (* ram_style = "distributed" *) reg [21:0] FetchCachePlugin_logic_ways_2_mem [0:63];
  (* ram_style = "distributed" *) reg [21:0] FetchCachePlugin_logic_ways_3_mem [0:63];
  (* ram_style = "distributed" *) reg [2:0] FetchCachePlugin_logic_plru_ram [0:63];
  (* ram_style = "distributed" *) reg [31:0] DecoderPredictionPlugin_logic_ras_mem_stack [0:15];
  reg [49:0] BtbPlugin_logic_mem [0:511];
  reg [3:0] GSharePlugin_logic_mem_counter [0:8191];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_lq_mem_addressPre [0:15];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_lq_mem_addressPost [0:15];
  (* ram_style = "distributed" *) reg [1:0] Lsu2Plugin_logic_lq_mem_size [0:15];
  (* ram_style = "distributed" *) reg [5:0] Lsu2Plugin_logic_lq_mem_physRd [0:15];
  (* ram_style = "distributed" *) reg [5:0] Lsu2Plugin_logic_lq_mem_robId [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_robIdMsb [0:15];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_lq_mem_pc [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_io [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_writeRd [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_lr [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_unsigned [0:15];
  reg [31:0] Lsu2Plugin_logic_lq_mem_data [0:15];
  reg [0:0] Lsu2Plugin_logic_lq_mem_spFpAddress [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_lq_mem_hazardPrediction_valid [0:15];
  (* ram_style = "distributed" *) reg [3:0] Lsu2Plugin_logic_lq_mem_hazardPrediction_delta [0:15];
  (* ram_style = "distributed" *) reg [2:0] Lsu2Plugin_logic_lq_mem_hazardPrediction_score [0:15];
  reg [5:0] Lsu2Plugin_logic_lq_mem_hitPrediction_counter [0:15];
  reg [22:0] Lsu2Plugin_logic_lq_hazardPrediction_mem [0:127];
  reg [5:0] Lsu2Plugin_logic_lq_hitPrediction_mem [0:1023];
  (* ram_style = "distributed" *) reg [5:0] Lsu2Plugin_logic_sq_mem_robId [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_robIdMsb [0:15];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_sq_mem_addressPre [0:15];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_sq_mem_addressPost [0:15];
  (* ram_style = "distributed" *) reg [1:0] Lsu2Plugin_logic_sq_mem_size [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_io [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_amo [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_sc [0:15];
  (* ram_style = "distributed" *) reg [31:0] Lsu2Plugin_logic_sq_mem_data [0:15];
  (* ram_style = "distributed" *) reg [0:0] Lsu2Plugin_logic_sq_mem_doNotBypass [0:15];
  (* ram_style = "distributed" *) reg [41:0] FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0 [0:31];
  (* ram_style = "distributed" *) reg [41:0] FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1 [0:31];
  (* ram_style = "distributed" *) reg [41:0] FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2 [0:31];
  (* ram_style = "distributed" *) reg [41:0] FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3 [0:31];
  (* ram_style = "distributed" *) reg [21:0] FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0 [0:31];
  (* ram_style = "distributed" *) reg [21:0] FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1 [0:31];
  (* ram_style = "distributed" *) reg [41:0] Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0 [0:31];
  (* ram_style = "distributed" *) reg [41:0] Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1 [0:31];
  (* ram_style = "distributed" *) reg [41:0] Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2 [0:31];
  (* ram_style = "distributed" *) reg [41:0] Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3 [0:31];
  (* ram_style = "distributed" *) reg [21:0] Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0 [0:31];
  (* ram_style = "distributed" *) reg [21:0] Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1 [0:31];
  (* ram_style = "distributed" *) reg [31:0] CsrRamPlugin_logic_mem [0:31];
  (* ram_style = "distributed" *) reg [1:0] RobPlugin_logic_completionMem_target [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_0 [0:63];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_1 [0:63];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_2 [0:63];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_3 [0:63];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_4 [0:63];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_5 [0:63];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_completionMem_hits_6 [0:63];
  (* ram_style = "distributed" *) reg [1:0] RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [31:0] RobPlugin_logic_storage_PC_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [31:0] RobPlugin_logic_storage_PC_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_WRITE_RD_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_WRITE_RD_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [11:0] RobPlugin_logic_storage_PHYS_RD_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [9:0] RobPlugin_logic_storage_ARCH_RD_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [11:0] RobPlugin_logic_storage_PHYS_RD_FREE_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [1:0] RobPlugin_logic_storage_BRANCH_SEL_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [23:0] RobPlugin_logic_storage_BRANCH_HISTORY_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [23:0] RobPlugin_logic_storage_BRANCH_HISTORY_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [3:0] RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [3:0] RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [1:0] RobPlugin_logic_storage_LQ_ALLOC_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [1:0] RobPlugin_logic_storage_SQ_ALLOC_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [31:0] RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [31:0] RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [5:0] RobPlugin_logic_storage_PHYS_RS_0_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [5:0] RobPlugin_logic_storage_PHYS_RS_0_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_READ_RS_0_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_READ_RS_0_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [5:0] RobPlugin_logic_storage_PHYS_RS_1_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [5:0] RobPlugin_logic_storage_PHYS_RS_1_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_READ_RS_1_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_READ_RS_1_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [3:0] RobPlugin_logic_storage_BRANCH_ID_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [3:0] RobPlugin_logic_storage_BRANCH_ID_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [4:0] RobPlugin_logic_storage_LSU_ID_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [4:0] RobPlugin_logic_storage_LSU_ID_banks_1 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_ROB_MSB_banks_0 [0:31];
  (* ram_style = "distributed" *) reg [0:0] RobPlugin_logic_storage_ROB_MSB_banks_1 [0:31];
  function [31:0] zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue(input dummy);
    begin
      zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue = 32'h00000000;
      zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue[2 : 0] = 3'b101;
    end
  endfunction
  wire [31:0] _zz_322;
  function  zz_DecoderPlugin_logic_slots_0_x0AlwaysZero(input dummy);
    begin
      zz_DecoderPlugin_logic_slots_0_x0AlwaysZero = 1'bx;
      zz_DecoderPlugin_logic_slots_0_x0AlwaysZero = 1'b1;
    end
  endfunction
  wire  _zz_323;
  function  zz_DecoderPlugin_logic_slots_1_x0AlwaysZero(input dummy);
    begin
      zz_DecoderPlugin_logic_slots_1_x0AlwaysZero = 1'bx;
      zz_DecoderPlugin_logic_slots_1_x0AlwaysZero = 1'b1;
    end
  endfunction
  wire  _zz_324;

  assign _zz_FetchPlugin_stages_1_FETCH_ID_1 = FetchPlugin_stages_1_isFireing;
  assign _zz_FetchPlugin_stages_1_FETCH_ID = {11'd0, _zz_FetchPlugin_stages_1_FETCH_ID_1};
  assign _zz_FetchCachePlugin_logic_refill_randomWay_valueNext_1 = FetchCachePlugin_logic_refill_randomWay_willIncrement;
  assign _zz_FetchCachePlugin_logic_refill_randomWay_valueNext = {1'd0, _zz_FetchCachePlugin_logic_refill_randomWay_valueNext_1};
  assign _zz_FetchCachePlugin_logic_read_onWays_0_hits_bypassHits = (FetchPlugin_stages_1_Fetch_FETCH_PC >>> 4'd12);
  assign _zz_FetchCachePlugin_logic_read_onWays_1_hits_bypassHits = (FetchPlugin_stages_1_Fetch_FETCH_PC >>> 4'd12);
  assign _zz_FetchCachePlugin_logic_read_onWays_2_hits_bypassHits = (FetchPlugin_stages_1_Fetch_FETCH_PC >>> 4'd12);
  assign _zz_FetchCachePlugin_logic_read_onWays_3_hits_bypassHits = (FetchPlugin_stages_1_Fetch_FETCH_PC >>> 4'd12);
  assign _zz_AlignerPlugin_logic_extractors_0_usable = (((_zz_AlignerPlugin_logic_extractors_0_usage ? AlignerPlugin_logic_decoders_0_usable : 1'b0) | (_zz_AlignerPlugin_logic_extractors_0_usage_1 ? AlignerPlugin_logic_decoders_1_usable : 1'b0)) | ((_zz_AlignerPlugin_logic_extractors_0_usage_2 ? AlignerPlugin_logic_decoders_2_usable : 1'b0) | (_zz_AlignerPlugin_logic_extractors_0_usage_3 ? AlignerPlugin_logic_decoders_3_usable : 1'b0)));
  assign _zz_FrontendPlugin_aligned_PC_0 = (AlignerPlugin_logic_extractors_0_pcWord >>> 2'd3);
  assign _zz_AlignerPlugin_logic_extractors_1_usable = (((_zz_AlignerPlugin_logic_extractors_1_usage ? AlignerPlugin_logic_decoders_1_usable : 1'b0) | (_zz_AlignerPlugin_logic_extractors_1_usage_1 ? AlignerPlugin_logic_decoders_2_usable : 1'b0)) | (_zz_AlignerPlugin_logic_extractors_1_usage_2 ? AlignerPlugin_logic_decoders_3_usable : 1'b0));
  assign _zz_FrontendPlugin_aligned_PC_1 = (AlignerPlugin_logic_extractors_1_pcWord >>> 2'd3);
  assign _zz_DispatchPlugin_logic_sparseRob_sparse_ohFirst_masked = (DispatchPlugin_logic_sparseRob_sparse_ohFirst_input - 2'b01);
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push = (DecoderPredictionPlugin_logic_ras_ptr_push + _zz_DecoderPredictionPlugin_logic_ras_ptr_push_1);
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push_2 = DecoderPredictionPlugin_logic_ras_ptr_pushIt;
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push_1 = {3'd0, _zz_DecoderPredictionPlugin_logic_ras_ptr_push_2};
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push_4 = DecoderPredictionPlugin_logic_ras_ptr_popIt;
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_push_3 = {3'd0, _zz_DecoderPredictionPlugin_logic_ras_ptr_push_4};
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop = (DecoderPredictionPlugin_logic_ras_ptr_pop + _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_1);
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_2 = DecoderPredictionPlugin_logic_ras_ptr_pushIt;
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_1 = {3'd0, _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_2};
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_4 = DecoderPredictionPlugin_logic_ras_ptr_popIt;
  assign _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_3 = {3'd0, _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_4};
  assign _zz_BtbPlugin_logic_onLearn_port_payload_address = (BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice >>> 2'd3);
  assign _zz_BtbPlugin_logic_onLearn_port_payload_data_slice = (BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice >>> 2'd2);
  assign _zz_BtbPlugin_logic_readCmd_entryAddress = (FetchPlugin_stages_0_Fetch_FETCH_PC >>> 2'd3);
  assign _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_5 = FetchPlugin_stages_0_BRANCH_HISTORY;
  assign _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_4 = _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_5[12:0];
  assign _zz_GSharePlugin_logic_onLearn_hash_5 = BranchContextPlugin_free_learn_BRANCH_HISTORY;
  assign _zz_GSharePlugin_logic_onLearn_hash_4 = _zz_GSharePlugin_logic_onLearn_hash_5[12:0];
  assign _zz_CommitPlugin_logic_ptr_allocNext_1 = (FrontendPlugin_allocated_isFireing ? 2'b10 : 2'b00);
  assign _zz_CommitPlugin_logic_ptr_allocNext = {5'd0, _zz_CommitPlugin_logic_ptr_allocNext_1};
  assign _zz_CommitPlugin_logic_reschedule_commit_rowHit = CommitPlugin_logic_ptr_commitRow[4:0];
  assign _zz_CommitPlugin_logic_reschedule_age = CommitPlugin_logic_ptr_free[5:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_0_age = CommitPlugin_logic_ptr_free[5:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_1_age = CommitPlugin_logic_ptr_free[5:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_2_age = CommitPlugin_logic_ptr_free[5:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_3_age = CommitPlugin_logic_ptr_free[5:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_4_age = CommitPlugin_logic_ptr_free[5:0];
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_5_age = CommitPlugin_logic_ptr_free[5:0];
  assign _zz_CommitPlugin_logic_reschedule_trap_6 = ((((_zz_CommitPlugin_logic_reschedule_trap ? Lsu2Plugin_setup_sharedTrap_payload_trap : 1'b0) | (_zz_CommitPlugin_logic_reschedule_trap_1 ? 1'b1 : 1'b0)) | ((_zz_CommitPlugin_logic_reschedule_trap_2 ? ALU0_BranchPlugin_setup_reschedule_payload_trap : 1'b0) | (_zz_CommitPlugin_logic_reschedule_trap_3 ? 1'b1 : 1'b0))) | ((_zz_CommitPlugin_logic_reschedule_trap_4 ? 1'b1 : 1'b0) | (_zz_CommitPlugin_logic_reschedule_trap_5 ? ALU1_BranchPlugin_setup_reschedule_payload_trap : 1'b0)));
  assign _zz_CommitPlugin_logic_reschedule_skipCommit = ((((CommitPlugin_logic_reschedule_portsLogic_hits[0] ? Lsu2Plugin_setup_sharedTrap_payload_skipCommit : 1'b0) | (CommitPlugin_logic_reschedule_portsLogic_hits[1] ? Lsu2Plugin_setup_specialTrap_payload_skipCommit : 1'b0)) | ((CommitPlugin_logic_reschedule_portsLogic_hits[2] ? ALU0_BranchPlugin_setup_reschedule_payload_skipCommit : 1'b0) | (CommitPlugin_logic_reschedule_portsLogic_hits[3] ? EnvCallPlugin_setup_reschedule_payload_skipCommit : 1'b0))) | ((CommitPlugin_logic_reschedule_portsLogic_hits[4] ? EU0_CsrAccessPlugin_setup_trap_payload_skipCommit : 1'b0) | (CommitPlugin_logic_reschedule_portsLogic_hits[5] ? ALU1_BranchPlugin_setup_reschedule_payload_skipCommit : 1'b0)));
  assign _zz__zz_CommitPlugin_logic_commit_head_1 = (_zz_CommitPlugin_logic_commit_head & (~ _zz__zz_CommitPlugin_logic_commit_head_1_1));
  assign _zz__zz_CommitPlugin_logic_commit_head_1_1 = (_zz_CommitPlugin_logic_commit_head - 2'b01);
  assign _zz_CommitPlugin_logic_commit_head_2 = (CommitPlugin_logic_ptr_commit + _zz_CommitPlugin_logic_commit_head_3);
  assign _zz_CommitPlugin_logic_commit_head_4 = _zz_CommitPlugin_logic_commit_head_1;
  assign _zz_CommitPlugin_logic_commit_head_3 = {6'd0, _zz_CommitPlugin_logic_commit_head_4};
  assign _zz_CommitPlugin_logic_free_robHit = CommitPlugin_logic_ptr_free[5:0];
  assign _zz_CommitDebugFilterPlugin_logic_filters_0_value = ($signed(_zz_CommitDebugFilterPlugin_logic_filters_0_value_1) >>> 4);
  assign _zz_CommitDebugFilterPlugin_logic_filters_0_value_1 = _zz_CommitDebugFilterPlugin_logic_filters_0_value_2;
  assign _zz_CommitDebugFilterPlugin_logic_filters_0_value_2 = (_zz_CommitDebugFilterPlugin_logic_filters_0_value_3 - CommitDebugFilterPlugin_logic_filters_0_value);
  assign _zz_CommitDebugFilterPlugin_logic_filters_0_value_3 = {14'd0, CommitDebugFilterPlugin_logic_commits};
  assign _zz_CommitDebugFilterPlugin_logic_filters_1_value = ($signed(_zz_CommitDebugFilterPlugin_logic_filters_1_value_1) >>> 8);
  assign _zz_CommitDebugFilterPlugin_logic_filters_1_value_1 = _zz_CommitDebugFilterPlugin_logic_filters_1_value_2;
  assign _zz_CommitDebugFilterPlugin_logic_filters_1_value_2 = (_zz_CommitDebugFilterPlugin_logic_filters_1_value_3 - CommitDebugFilterPlugin_logic_filters_1_value);
  assign _zz_CommitDebugFilterPlugin_logic_filters_1_value_3 = {14'd0, CommitDebugFilterPlugin_logic_commits};
  assign _zz_CommitDebugFilterPlugin_logic_filters_2_value = ($signed(_zz_CommitDebugFilterPlugin_logic_filters_2_value_1) >>> 12);
  assign _zz_CommitDebugFilterPlugin_logic_filters_2_value_1 = _zz_CommitDebugFilterPlugin_logic_filters_2_value_2;
  assign _zz_CommitDebugFilterPlugin_logic_filters_2_value_2 = (_zz_CommitDebugFilterPlugin_logic_filters_2_value_3 - CommitDebugFilterPlugin_logic_filters_2_value);
  assign _zz_CommitDebugFilterPlugin_logic_filters_2_value_3 = {14'd0, CommitDebugFilterPlugin_logic_commits};
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2 = {4'd0, PerformanceCounterPlugin_logic_commitCount_regNext};
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3_1 = ((((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_7 == 3'b001) ? PerformanceCounterPlugin_logic_events_sums_0 : 1'b0) | ((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_7 == 3'b010) ? PerformanceCounterPlugin_logic_events_sums_1 : 1'b0)) | (((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_7 == 3'b011) ? PerformanceCounterPlugin_logic_events_sums_2 : 1'b0) | ((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_7 == 3'b100) ? PerformanceCounterPlugin_logic_events_sums_3 : 1'b0)));
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3 = {5'd0, _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3_1};
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4_1 = ((((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_8 == 3'b001) ? PerformanceCounterPlugin_logic_events_sums_0 : 1'b0) | ((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_8 == 3'b010) ? PerformanceCounterPlugin_logic_events_sums_1 : 1'b0)) | (((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_8 == 3'b011) ? PerformanceCounterPlugin_logic_events_sums_2 : 1'b0) | ((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_8 == 3'b100) ? PerformanceCounterPlugin_logic_events_sums_3 : 1'b0)));
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4 = {5'd0, _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4_1};
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5_1 = ((((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_9 == 3'b001) ? PerformanceCounterPlugin_logic_events_sums_0 : 1'b0) | ((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_9 == 3'b010) ? PerformanceCounterPlugin_logic_events_sums_1 : 1'b0)) | (((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_9 == 3'b011) ? PerformanceCounterPlugin_logic_events_sums_2 : 1'b0) | ((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_9 == 3'b100) ? PerformanceCounterPlugin_logic_events_sums_3 : 1'b0)));
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5 = {5'd0, _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5_1};
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6_1 = ((((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_10 == 3'b001) ? PerformanceCounterPlugin_logic_events_sums_0 : 1'b0) | ((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_10 == 3'b010) ? PerformanceCounterPlugin_logic_events_sums_1 : 1'b0)) | (((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_10 == 3'b011) ? PerformanceCounterPlugin_logic_events_sums_2 : 1'b0) | ((_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_10 == 3'b100) ? PerformanceCounterPlugin_logic_events_sums_3 : 1'b0)));
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6 = {5'd0, _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6_1};
  assign _zz__zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1) + $signed(ALU0_SrcPlugin_logic_addsub_rs2Patched));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1 = _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2 = {31'd0, _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3};
  assign _zz_ALU0_IntAluPlugin_logic_process_result_1 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
  assign _zz_ALU0_IntAluPlugin_logic_process_result = {31'd0, _zz_ALU0_IntAluPlugin_logic_process_result_1};
  assign _zz_ALU0_ShiftPlugin_logic_process_amplitude = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[4 : 0];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed = {ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[0],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[1],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[2],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[3],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[4],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[5],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[6],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[7],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[8],{_zz_ALU0_ShiftPlugin_logic_process_reversed_1,{_zz_ALU0_ShiftPlugin_logic_process_reversed_2,_zz_ALU0_ShiftPlugin_logic_process_reversed_3}}}}}}}}}}};
  assign _zz_ALU0_ShiftPlugin_logic_process_shifted = ($signed(_zz_ALU0_ShiftPlugin_logic_process_shifted_1) >>> ALU0_ShiftPlugin_logic_process_amplitude);
  assign _zz_ALU0_ShiftPlugin_logic_process_shifted_1 = {(ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SIGNED && ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]),ALU0_ShiftPlugin_logic_process_reversed};
  assign _zz_ALU0_ShiftPlugin_logic_process_patched = {ALU0_ShiftPlugin_logic_process_shifted[0],{ALU0_ShiftPlugin_logic_process_shifted[1],{ALU0_ShiftPlugin_logic_process_shifted[2],{ALU0_ShiftPlugin_logic_process_shifted[3],{ALU0_ShiftPlugin_logic_process_shifted[4],{ALU0_ShiftPlugin_logic_process_shifted[5],{ALU0_ShiftPlugin_logic_process_shifted[6],{ALU0_ShiftPlugin_logic_process_shifted[7],{ALU0_ShiftPlugin_logic_process_shifted[8],{_zz_ALU0_ShiftPlugin_logic_process_patched_1,{_zz_ALU0_ShiftPlugin_logic_process_patched_2,_zz_ALU0_ShiftPlugin_logic_process_patched_3}}}}}}}}}}};
  assign _zz_ALU0_BranchPlugin_logic_process_target_b = {{{{ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31],ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[19 : 12]},ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[20]},ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[30 : 21]},1'b0};
  assign _zz_ALU0_BranchPlugin_logic_process_target_b_1 = ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_ALU0_BranchPlugin_logic_process_target_b_2 = {{{{ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31],ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[7]},ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[30 : 25]},ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[11 : 8]},1'b0};
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE = ($signed(ALU0_BranchPlugin_logic_process_target_a) + $signed(ALU0_BranchPlugin_logic_process_target_b));
  assign _zz_ALU0_BranchPlugin_logic_process_slices_1 = 1'b0;
  assign _zz_ALU0_BranchPlugin_logic_process_slices = {1'd0, _zz_ALU0_BranchPlugin_logic_process_slices_1};
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE_1 = ({2'd0,ALU0_BranchPlugin_logic_process_slices} <<< 2'd2);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE = {28'd0, _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE_1};
  assign _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = {EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 25],EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[11 : 7]};
  assign _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2_1 = EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1) + $signed(EU0_SrcPlugin_logic_addsub_rs2Patched));
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3 = EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2 = {31'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED_1 = EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED = {31'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED_1 = EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED = {31'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_1 = ($signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_2) * $signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_3));
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1 = {{13{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_1[33]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_2 = {1'b0,EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[16 : 0]};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1_3 = EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[32 : 17];
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_1 = ($signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_2) * $signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_3));
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2 = {{13{_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_1[33]}}, _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_2 = EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 17];
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2_3 = {1'b0,EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[16 : 0]};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3_1 = ($signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3_2) * $signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3_3));
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3_1[29:0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3_2 = EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[32 : 17];
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3_3 = EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[32 : 17];
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_3 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_5);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_4 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_2};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_3 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_4 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_5);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_4 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_5 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_1};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_6 = {2'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_2};
  assign _zz_EU0_DivPlugin_logic_rsp_selected = {2'd0, EU0_DivPlugin_logic_div_io_rsp_payload_remain};
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_1 = _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_2;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_2 = ((EU0_ExecutionUnitBase_pipeline_execute_1_DIV_REVERT_RESULT ? (~ _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT) : _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT) + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_3);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_4 = EU0_ExecutionUnitBase_pipeline_execute_1_DIV_REVERT_RESULT;
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_3 = {34'd0, _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_4};
  assign _zz__zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1) + $signed(ALU1_SrcPlugin_logic_addsub_rs2Patched));
  assign _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1 = _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2;
  assign _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3 = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT;
  assign _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_2 = {31'd0, _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_3};
  assign _zz_ALU1_IntAluPlugin_logic_process_result_1 = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
  assign _zz_ALU1_IntAluPlugin_logic_process_result = {31'd0, _zz_ALU1_IntAluPlugin_logic_process_result_1};
  assign _zz_ALU1_ShiftPlugin_logic_process_amplitude = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[4 : 0];
  assign _zz_ALU1_ShiftPlugin_logic_process_reversed = {ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[0],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[1],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[2],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[3],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[4],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[5],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[6],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[7],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[8],{_zz_ALU1_ShiftPlugin_logic_process_reversed_1,{_zz_ALU1_ShiftPlugin_logic_process_reversed_2,_zz_ALU1_ShiftPlugin_logic_process_reversed_3}}}}}}}}}}};
  assign _zz_ALU1_ShiftPlugin_logic_process_shifted = ($signed(_zz_ALU1_ShiftPlugin_logic_process_shifted_1) >>> ALU1_ShiftPlugin_logic_process_amplitude);
  assign _zz_ALU1_ShiftPlugin_logic_process_shifted_1 = {(ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SIGNED && ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]),ALU1_ShiftPlugin_logic_process_reversed};
  assign _zz_ALU1_ShiftPlugin_logic_process_patched = {ALU1_ShiftPlugin_logic_process_shifted[0],{ALU1_ShiftPlugin_logic_process_shifted[1],{ALU1_ShiftPlugin_logic_process_shifted[2],{ALU1_ShiftPlugin_logic_process_shifted[3],{ALU1_ShiftPlugin_logic_process_shifted[4],{ALU1_ShiftPlugin_logic_process_shifted[5],{ALU1_ShiftPlugin_logic_process_shifted[6],{ALU1_ShiftPlugin_logic_process_shifted[7],{ALU1_ShiftPlugin_logic_process_shifted[8],{_zz_ALU1_ShiftPlugin_logic_process_patched_1,{_zz_ALU1_ShiftPlugin_logic_process_patched_2,_zz_ALU1_ShiftPlugin_logic_process_patched_3}}}}}}}}}}};
  assign _zz_ALU1_BranchPlugin_logic_process_target_b = {{{{ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31],ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[19 : 12]},ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[20]},ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[30 : 21]},1'b0};
  assign _zz_ALU1_BranchPlugin_logic_process_target_b_1 = ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_ALU1_BranchPlugin_logic_process_target_b_2 = {{{{ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31],ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[7]},ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[30 : 25]},ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[11 : 8]},1'b0};
  assign _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TRUE = ($signed(ALU1_BranchPlugin_logic_process_target_a) + $signed(ALU1_BranchPlugin_logic_process_target_b));
  assign _zz_ALU1_BranchPlugin_logic_process_slices_1 = 1'b0;
  assign _zz_ALU1_BranchPlugin_logic_process_slices = {1'd0, _zz_ALU1_BranchPlugin_logic_process_slices_1};
  assign _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE_1 = ({2'd0,ALU1_BranchPlugin_logic_process_slices} <<< 2'd2);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE = {28'd0, _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE_1};
  assign _zz_BranchContextPlugin_logic_onCommit_commitedNext = {3'd0, _zz_BranchContextPlugin_logic_onCommit_commitedNext_1};
  assign _zz_HistoryPlugin_logic_onCommit_valueNext_1 = {HistoryPlugin_logic_onCommit_valueNext,HistoryPlugin_logic_onCommit_isTaken_0};
  assign _zz_HistoryPlugin_logic_onCommit_valueNext_2 = {HistoryPlugin_logic_onCommit_valueNext_1,HistoryPlugin_logic_onCommit_isTaken_1};
  assign _zz_HistoryPlugin_logic_update_pushes_0_stateNext_1 = {HistoryPlugin_logic_update_pushes_0_stateNext,BtbPlugin_setup_historyPush_taken[0]};
  assign _zz_HistoryPlugin_logic_update_pushes_2_stateNext_1 = {HistoryPlugin_logic_update_pushes_2_stateNext,DecoderPredictionPlugin_setup_historyPush_taken[0]};
  assign _zz_HistoryPlugin_logic_update_pushes_2_stateNext_2 = {HistoryPlugin_logic_update_pushes_2_stateNext_1,DecoderPredictionPlugin_setup_historyPush_taken[1]};
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken = _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken_1[0 : 0];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken_1 = RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_2_rsp[0];
  assign _zz_Lsu2Plugin_logic_lq_tracker_freeNext = (Lsu2Plugin_logic_lq_tracker_free + _zz_Lsu2Plugin_logic_lq_tracker_freeNext_1);
  assign _zz_Lsu2Plugin_logic_lq_tracker_freeNext_1 = {3'd0, Lsu2Plugin_logic_lq_tracker_add};
  assign _zz_Lsu2Plugin_logic_lq_tracker_freeNext_2 = {3'd0, Lsu2Plugin_logic_lq_tracker_sub};
  assign _zz_when_Lsu2Plugin_l454 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_1 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_2 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_3 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_4 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_5 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_6 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_7 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_8 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_9 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_10 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_11 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_12 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_13 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_14 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_when_Lsu2Plugin_l454_15 = Lsu2Plugin_logic_lq_onCommit_free[3:0];
  assign _zz_Lsu2Plugin_logic_lq_onCommit_priority_1 = (Lsu2Plugin_logic_lq_onCommit_priority <<< 1);
  assign _zz_Lsu2Plugin_logic_lq_onCommit_free_1_1 = Lsu2Plugin_logic_lq_onCommit_lqCommits_0;
  assign _zz_Lsu2Plugin_logic_lq_onCommit_free_1 = {4'd0, _zz_Lsu2Plugin_logic_lq_onCommit_free_1_1};
  assign _zz_when_Lsu2Plugin_l454_16 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_17 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_18 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_19 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_20 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_21 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_22 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_23 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_24 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_25 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_26 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_27 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_28 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_29 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_30 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_when_Lsu2Plugin_l454_31 = Lsu2Plugin_logic_lq_onCommit_free_1[3:0];
  assign _zz_Lsu2Plugin_logic_lq_onCommit_priority_2 = (Lsu2Plugin_logic_lq_onCommit_priority_1 <<< 1);
  assign _zz_Lsu2Plugin_logic_lq_onCommit_free_2_1 = Lsu2Plugin_logic_lq_onCommit_lqCommits_1;
  assign _zz_Lsu2Plugin_logic_lq_onCommit_free_2 = {4'd0, _zz_Lsu2Plugin_logic_lq_onCommit_free_2_1};
  assign _zz_Lsu2Plugin_logic_lq_ptr_free = {3'd0, Lsu2Plugin_logic_lq_onCommit_lqCommitCount};
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext = (_zz_Lsu2Plugin_logic_sq_tracker_freeNext_1 - _zz_Lsu2Plugin_logic_sq_tracker_freeNext_3);
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext_1 = (_zz_Lsu2Plugin_logic_sq_tracker_freeNext_2 - Lsu2Plugin_logic_sq_ptr_alloc);
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext_2 = (5'h10 + Lsu2Plugin_logic_sq_ptr_free);
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext_3 = {3'd0, Lsu2Plugin_logic_sq_tracker_sub};
  assign _zz_Lsu2Plugin_logic_sq_tracker_freeNext_4 = {4'd0, Lsu2Plugin_logic_sq_tracker_add};
  assign _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1_1 = when_Lsu2Plugin_l591;
  assign _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1 = {4'd0, _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1_1};
  assign _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_2_1 = when_Lsu2Plugin_l591_1;
  assign _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_2 = {4'd0, _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_2_1};
  assign _zz_Lsu2Plugin_logic_lq_mem_addressPre_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_physRd_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_robId_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_pc_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_writeRd_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_lr_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_size_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_unsigned_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_addressPre_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_robId_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_amo_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_sc_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_size_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_data_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh = ({1'd0,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pHigh} <<< 1'd1);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh = ({1'd0,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pHigh} <<< 1'd1);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s1_cmp = (Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ROB_FULL - Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ROB_FULL);
  assign _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu = ({AguPlugin_setup_port_payload_robIdMsb,AguPlugin_setup_port_payload_robId} - Lsu2Plugin_logic_sharedPip_stages_0_LQ_ROB_FULL);
  assign _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu_1 = ({AguPlugin_setup_port_payload_robIdMsb,AguPlugin_setup_port_payload_robId} - Lsu2Plugin_logic_sharedPip_stages_0_SQ_ROB_FULL);
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID = ((Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ || (! Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask)) ? Lsu2Plugin_logic_sharedPip_stages_0_LQ_ROB_FULL : Lsu2Plugin_logic_sharedPip_stages_0_SQ_ROB_FULL);
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_1 = {AguPlugin_setup_port_payload_robIdMsb,AguPlugin_setup_port_payload_robId};
  assign _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT = (Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC - _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1);
  assign _zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1 = {1'd0, Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA};
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1 = (_zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT - Lsu2Plugin_logic_sq_ptr_free);
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh = {1'd0, Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pLow};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh = ({1'd0,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pHigh} <<< 1'd1);
  assign _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta = (_zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_1 - 5'h01);
  assign _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_1 = (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_3_rsp - _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_2);
  assign _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta_2 = {1'd0, Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID};
  assign _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_1 = {Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION_COUNTER[5],Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION_COUNTER};
  assign _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_2 = {_zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[5],_zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next};
  assign _zz_when_SInt_l132 = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[6 : 5];
  assign _zz_when_SInt_l138 = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[5 : 5];
  assign _zz_Lsu2Plugin_logic_sq_ptr_writeBack_1 = Lsu2Plugin_logic_writeback_feed_fire;
  assign _zz_Lsu2Plugin_logic_sq_ptr_writeBack = {4'd0, _zz_Lsu2Plugin_logic_sq_ptr_writeBack_1};
  assign _zz_Lsu2Plugin_setup_specialTrap_payload_cause = (Lsu2Plugin_logic_special_isStore ? 3'b111 : 3'b101);
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_2 = ($signed(_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_3) + $signed(_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_6));
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_3 = ($signed(_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_4) + $signed(_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_5));
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_4 = _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1;
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_5 = (Lsu2Plugin_logic_special_atomic_alu_compare ? (~ _zz_Lsu2Plugin_logic_special_atomic_alu_addSub) : _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_7 = (Lsu2Plugin_logic_special_atomic_alu_compare ? 2'b01 : 2'b00);
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_6 = {{30{_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_7[1]}}, _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_7};
  assign _zz_ALU0_BranchPlugin_setup_intFormatPort_payload = ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE;
  assign _zz_ALU0_BranchPlugin_setup_reschedule_payload_reason = ((ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL == BranchPlugin_BranchCtrlEnum_B) ? 5'h10 : 5'h11);
  assign _zz_ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice_1 = 2'b00;
  assign _zz_ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice = {30'd0, _zz_ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice_1};
  assign _zz_ALU1_BranchPlugin_setup_intFormatPort_payload = ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE;
  assign _zz_ALU1_BranchPlugin_setup_reschedule_payload_reason = ((ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL == BranchPlugin_BranchCtrlEnum_B) ? 5'h10 : 5'h11);
  assign _zz_ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice_1 = 2'b00;
  assign _zz_ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice = {30'd0, _zz_ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice_1};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement;
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext = {1'd0, _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement;
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext = {1'd0, _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext_1};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_6 = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowExecute : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowExecute : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowExecute : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowExecute : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowExecute : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowExecute : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowRead : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowRead : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowRead : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowRead : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowRead : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowRead : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowWrite : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowWrite : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowWrite : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowWrite : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowWrite : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowWrite : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowUser : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowUser : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowUser : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowUser : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowUser : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowUser : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_pageFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_pageFault : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_pageFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_pageFault : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_pageFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_pageFault : 1'b0)));
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_accessFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_accessFault : 1'b0)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_accessFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_accessFault : 1'b0))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_accessFault : 1'b0) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_accessFault : 1'b0)));
  assign _zz_PerformanceCounterPlugin_setup_readPort_address = {2'd0, PerformanceCounterPlugin_logic_fsm_cmd_address};
  assign _zz_PerformanceCounterPlugin_setup_writePort_address = {2'd0, PerformanceCounterPlugin_logic_fsm_cmd_address};
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc = (PerformanceCounterPlugin_logic_fsm_ramReaded[63 : 5] + _zz_PerformanceCounterPlugin_logic_fsm_calc_1);
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_2 = PerformanceCounterPlugin_logic_fsm_counterReaded[5];
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_1 = {58'd0, _zz_PerformanceCounterPlugin_logic_fsm_calc_2};
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_3 = PerformanceCounterPlugin_logic_fsm_counterReaded[4:0];
  assign _zz_PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked = (PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input - 7'h01);
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_6 = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowExecute : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowExecute : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowExecute : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowExecute : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowExecute : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowExecute : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowRead : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowRead : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowRead : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowRead : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowRead : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowRead : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowWrite : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowWrite : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowWrite : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowWrite : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowWrite : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowWrite : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowUser : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowUser : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowUser : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowUser : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowUser : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowUser : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineException = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_pageFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_pageFault : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_pageFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_pageFault : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_pageFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_pageFault : 1'b0)));
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? FetchPlugin_stages_1_MMU_L0_ENTRIES_0_accessFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_1_accessFault : 1'b0)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_2_accessFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? FetchPlugin_stages_1_MMU_L0_ENTRIES_3_accessFault : 1'b0))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_0_accessFault : 1'b0) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? FetchPlugin_stages_1_MMU_L1_ENTRIES_1_accessFault : 1'b0)));
  assign _zz_MmuPlugin_logic_refill_portsRequests_ohFirst_masked = (MmuPlugin_logic_refill_portsRequests_ohFirst_input - 2'b01);
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask_1 = (4'b0001 <<< FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value);
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask_1 = (4'b0001 <<< Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value);
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask = (2'b01 <<< FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value);
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask = (2'b01 <<< Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value);
  assign _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input - 4'b0001);
  assign _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input - 3'b001);
  assign _zz_EU0_CsrAccessPlugin_setup_onDecodeAddress = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
  assign _zz_EU0_CsrAccessPlugin_setup_onReadAddress = EU0_CsrAccessPlugin_logic_fsm_regs_microOp;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1 = EU0_CsrAccessPlugin_logic_fsm_regs_microOp[19 : 15];
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = {27'd0, _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1};
  assign _zz_EU0_CsrAccessPlugin_setup_onWriteAddress = EU0_CsrAccessPlugin_logic_fsm_regs_microOp;
  assign _zz_csrAccess_payload_address = EU0_ExecutionUnitBase_pipeline_execute_2_Frontend_MICRO_OP;
  assign _zz_FrontendPlugin_decoded_READ_RS_0_0 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000044) == 32'h00000000),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000018) == 32'h00000000),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00006004) == 32'h00002000),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00005004) == 32'h00001000),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00002050) == 32'h00002000)}}}});
  assign _zz_FrontendPlugin_decoded_READ_RS_1_0 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000034) == 32'h00000020),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000064) == 32'h00000020),{_zz_FrontendPlugin_decoded_SQ_ALLOC_0_1,_zz_FrontendPlugin_decoded_SQ_ALLOC_0}}});
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_1 = (|{_zz_FrontendPlugin_decoded_WRITE_RD_0,{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00001010) == 32'h00001010),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00002010) == 32'h00002010),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_WRITE_RD_0_2) == 32'h00002008),{(_zz_FrontendPlugin_decoded_WRITE_RD_0_3 == _zz_FrontendPlugin_decoded_WRITE_RD_0_4),{_zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_0,_zz_FrontendPlugin_decoded_WRITE_RD_0_5}}}}}});
  assign _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_0_1 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000030) == 32'h00000010),{_zz_FrontendPlugin_decoded_IS_ANY_0,{_zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_0,((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h02000050) == 32'h00000010)}}});
  assign _zz_FrontendPlugin_decoded_EU0_SEL_0 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000050) == 32'h00000050),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000050) == 32'h00000000),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h02000064) == 32'h02000020)}});
  assign _zz_FrontendPlugin_decoded_LQ_ALLOC_0 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000038) == 32'h00000000),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h18002048) == 32'h10002008)});
  assign _zz_FrontendPlugin_decoded_SQ_ALLOC_0_2 = (|{_zz_FrontendPlugin_decoded_SQ_ALLOC_0_1,{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000078) == 32'h00000020),_zz_FrontendPlugin_decoded_SQ_ALLOC_0}});
  assign _zz_FrontendPlugin_decoded_READ_RS_0_1 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000044) == 32'h00000000),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000018) == 32'h00000000),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00006004) == 32'h00002000),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00005004) == 32'h00001000),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00002050) == 32'h00002000)}}}});
  assign _zz_FrontendPlugin_decoded_READ_RS_1_1 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000034) == 32'h00000020),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000064) == 32'h00000020),{_zz_FrontendPlugin_decoded_SQ_ALLOC_1_1,_zz_FrontendPlugin_decoded_SQ_ALLOC_1}}});
  assign _zz_FrontendPlugin_decoded_WRITE_RD_1 = (|{_zz_FrontendPlugin_decoded_IS_JAL_1,{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00001010) == 32'h00001010),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00002010) == 32'h00002010),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & _zz_FrontendPlugin_decoded_WRITE_RD_1_1) == 32'h00002008),{(_zz_FrontendPlugin_decoded_WRITE_RD_1_2 == _zz_FrontendPlugin_decoded_WRITE_RD_1_3),{_zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_1,_zz_FrontendPlugin_decoded_WRITE_RD_1_4}}}}}});
  assign _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_1_1 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000030) == 32'h00000010),{_zz_FrontendPlugin_decoded_IS_ANY_1,{_zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_1,((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h02000050) == 32'h00000010)}}});
  assign _zz_FrontendPlugin_decoded_EU0_SEL_1 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000050) == 32'h00000050),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000050) == 32'h00000000),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h02000064) == 32'h02000020)}});
  assign _zz_FrontendPlugin_decoded_LQ_ALLOC_1 = (|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000038) == 32'h00000000),((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h18002048) == 32'h10002008)});
  assign _zz_FrontendPlugin_decoded_SQ_ALLOC_1_2 = (|{_zz_FrontendPlugin_decoded_SQ_ALLOC_1_1,{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000078) == 32'h00000020),_zz_FrontendPlugin_decoded_SQ_ALLOC_1}});
  assign _zz__zz_DecoderPlugin_setup_exceptionPort_payload_tval_1 = (_zz_DecoderPlugin_setup_exceptionPort_payload_tval & (~ _zz__zz_DecoderPlugin_setup_exceptionPort_payload_tval_1_1));
  assign _zz__zz_DecoderPlugin_setup_exceptionPort_payload_tval_1_1 = (_zz_DecoderPlugin_setup_exceptionPort_payload_tval - 2'b01);
  assign _zz_DecoderPlugin_logic_exception_fetchFault = ((DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_fetchFaultReg_0 : 1'b0) | (_zz_DecoderPlugin_setup_exceptionPort_payload_tval_1 ? DecoderPlugin_logic_exception_fetchFaultReg_1 : 1'b0));
  assign _zz_DecoderPlugin_logic_exception_fetchFaultPage = ((DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_fetchFaultPageReg_0 : 1'b0) | (_zz_DecoderPlugin_setup_exceptionPort_payload_tval_1 ? DecoderPlugin_logic_exception_fetchFaultPageReg_1 : 1'b0));
  assign _zz_DecoderPlugin_logic_exception_debugEnter = ((DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_debugEnterReg_0 : 1'b0) | (_zz_DecoderPlugin_setup_exceptionPort_payload_tval_1 ? DecoderPlugin_logic_exception_debugEnterReg_1 : 1'b0));
  assign _zz_DecoderPlugin_setup_exceptionPort_payload_tval_2 = (DecoderPlugin_logic_exception_pc + _zz_DecoderPlugin_setup_exceptionPort_payload_tval_3);
  assign _zz_DecoderPlugin_setup_exceptionPort_payload_tval_4 = 2'b00;
  assign _zz_DecoderPlugin_setup_exceptionPort_payload_tval_3 = {30'd0, _zz_DecoderPlugin_setup_exceptionPort_payload_tval_4};
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_2 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_3[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_3 = (|{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0,((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h10002048) == 32'h10002008)}}}});
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_2 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_3[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_3 = (|{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0,{((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h08002048) == 32'h08002008),((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h10002048) == 32'h00002008)}}});
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0 = _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_1[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0_1 = (|{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0,{((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h00002048) == 32'h00002008),_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0}}}});
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0_1[0];
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0_1 = 1'b0;
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0_1[0];
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0_1 = 1'b0;
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_2 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_3[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_3 = (|{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1,((FrontendPlugin_serialized_Frontend_MICRO_OP_1 & 32'h10002048) == 32'h10002008)}}}});
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_2 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_3[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_3 = (|{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1,{((FrontendPlugin_serialized_Frontend_MICRO_OP_1 & 32'h08002048) == 32'h08002008),((FrontendPlugin_serialized_Frontend_MICRO_OP_1 & 32'h10002048) == 32'h00002008)}}});
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_1 = _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_1_1[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_1_1 = (|{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_1,{_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1,{((FrontendPlugin_serialized_Frontend_MICRO_OP_1 & 32'h00002048) == 32'h00002008),_zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1}}}});
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_1 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_1_1[0];
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_1_1 = 1'b0;
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_1 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_1_1[0];
  assign _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_1_1 = 1'b0;
  assign _zz_FrontendPlugin_decoded_OP_ID_1 = ({1'd0,FrontendPlugin_decoded_isFireing} <<< 1'd1);
  assign _zz_FrontendPlugin_decoded_OP_ID = {10'd0, _zz_FrontendPlugin_decoded_OP_ID_1};
  assign _zz_FrontendPlugin_decoded_IS_JAL_0 = (|_zz_FrontendPlugin_decoded_WRITE_RD_0);
  assign _zz_FrontendPlugin_decoded_IS_JALR_0 = (|((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000001c) == 32'h00000004));
  assign _zz_FrontendPlugin_decoded_Prediction_IS_BRANCH_0 = (|((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000054) == 32'h00000040));
  assign _zz_FrontendPlugin_decoded_IS_ANY_0_1 = (|_zz_FrontendPlugin_decoded_IS_ANY_0);
  assign _zz__zz_FrontendPlugin_decoded_OFFSET_0 = {{{{FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[31],FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[7]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[30 : 25]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[11 : 8]},1'b0};
  assign _zz__zz_FrontendPlugin_decoded_OFFSET_0_1 = {{{{FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[31],FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[19 : 12]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[20]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[30 : 21]},1'b0};
  assign _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices_1 = 1'b0;
  assign _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices = {1'd0, _zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices_1};
  assign _zz_FrontendPlugin_decoded_PC_INC_0 = (FrontendPlugin_decoded_PC_0 + _zz_FrontendPlugin_decoded_PC_INC_0_1);
  assign _zz_FrontendPlugin_decoded_PC_INC_0_2 = ({2'd0,DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices} <<< 2'd2);
  assign _zz_FrontendPlugin_decoded_PC_INC_0_1 = {28'd0, _zz_FrontendPlugin_decoded_PC_INC_0_2};
  assign _zz_FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0 = FrontendPlugin_decoded_PC_0;
  assign _zz_FrontendPlugin_decoded_IS_JAL_1_1 = (|_zz_FrontendPlugin_decoded_IS_JAL_1);
  assign _zz_FrontendPlugin_decoded_IS_JALR_1 = (|((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000001c) == 32'h00000004));
  assign _zz_FrontendPlugin_decoded_Prediction_IS_BRANCH_1 = (|((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000054) == 32'h00000040));
  assign _zz_FrontendPlugin_decoded_IS_ANY_1_1 = (|_zz_FrontendPlugin_decoded_IS_ANY_1);
  assign _zz__zz_FrontendPlugin_decoded_OFFSET_1 = {{{{FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[31],FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[7]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[30 : 25]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[11 : 8]},1'b0};
  assign _zz__zz_FrontendPlugin_decoded_OFFSET_1_1 = {{{{FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[31],FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[19 : 12]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[20]},FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[30 : 21]},1'b0};
  assign _zz_DecoderPredictionPlugin_logic_decodePatch_slots_1_pcAdd_slices_1 = 1'b0;
  assign _zz_DecoderPredictionPlugin_logic_decodePatch_slots_1_pcAdd_slices = {1'd0, _zz_DecoderPredictionPlugin_logic_decodePatch_slots_1_pcAdd_slices_1};
  assign _zz_FrontendPlugin_decoded_PC_INC_1 = (FrontendPlugin_decoded_PC_1 + _zz_FrontendPlugin_decoded_PC_INC_1_1);
  assign _zz_FrontendPlugin_decoded_PC_INC_1_2 = ({2'd0,DecoderPredictionPlugin_logic_decodePatch_slots_1_pcAdd_slices} <<< 2'd2);
  assign _zz_FrontendPlugin_decoded_PC_INC_1_1 = {28'd0, _zz_FrontendPlugin_decoded_PC_INC_1_2};
  assign _zz_FrontendPlugin_decoded_PC_TARGET_PRE_RAS_1 = FrontendPlugin_decoded_PC_1;
  assign _zz_DecoderPredictionPlugin_setup_decodeJump_payload_pc = (FrontendPlugin_serialized_NEED_CORRECTION_0 ? FrontendPlugin_serialized_PC_PREDICTION_0 : FrontendPlugin_serialized_PC_PREDICTION_1);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2[31 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2 = _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port1[31 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_2[5 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_2 = _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port1[5 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2[0 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2 = _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_2[5 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_2 = _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port1[5 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2[0 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2 = _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2[0 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2 = _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port3[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_2[31 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_2 = _zz_RobPlugin_logic_storage_PC_banks_0_port3[31 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_2[3 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_2 = _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port1[3 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_2[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_2 = (|{((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002040) == 32'h00002000),{_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL,((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001040) == 32'h00000000)}});
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000040) == 32'h00000000));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00003044) == 32'h00001000));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004000) == 32'h00000000));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h40000000) == 32'h40000000));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL_1 = (|_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1_1 = (|_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_2[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_2 = (|{_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT,{((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002004) == 32'h00002000),((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h40000024) == 32'h40000020)}});
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1 = (|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000024) == 32'h00000024));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1 = (|{((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002010) == 32'h00002000),((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00005000) == 32'h00001000)});
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2[31 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2 = _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1_port1[31 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_2[5 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_2 = _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_1_port1[5 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2[0 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2 = _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_2[5 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_2 = _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_1_port1[5 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2[0 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2 = _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2[0 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2 = _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port3[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PC_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PC_2[31 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PC_2 = _zz_RobPlugin_logic_storage_PC_banks_1_port3[31 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_2[3 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_2 = _zz_RobPlugin_logic_storage_BRANCH_ID_banks_1_port1[3 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_2[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_2 = (|{((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002040) == 32'h00002000),{_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL,((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001040) == 32'h00000000)}});
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0_1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0_1 = (|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000040) == 32'h00000000));
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL_1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL_1 = (|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00003044) == 32'h00001000));
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT_1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT_1 = (|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004000) == 32'h00000000));
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED_1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED_1 = (|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h40000000) == 32'h40000000));
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL_1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL_1 = (|_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1_1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1_1 = (|_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_2[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_2 = (|{_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT,{((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002004) == 32'h00002000),((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h40000024) == 32'h40000020)}});
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1 = (|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000024) == 32'h00000024));
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED_1 = (|{((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002010) == 32'h00002000),((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00005000) == 32'h00001000)});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004050) == 32'h00000010));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2_1 = (|{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000010) == 32'h00000010),((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002008) == 32'h00000008)});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH_1 = (|{_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR,_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED_1 = (|{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001000) == 32'h00000000),_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_2 = (|{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00005000) == 32'h00004000),_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004060) == 32'h00004020));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM_1 = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL_1 = (|{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002010) == 32'h00002000),((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000018) == 32'h00000000)});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h10000008) == 32'h00000008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h10000008) == 32'h10000008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_2 = (|{_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD,((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h18000008) == 32'h10000008)});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT_1 = 1'b0;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000020) == 32'h00000020));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h10103040) == 32'h00000040));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h10103040) == 32'h00100040));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h12403040) == 32'h10000040));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h12203040) == 32'h10000040));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00003008) == 32'h00000008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00005008) == 32'h00001008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h02003040) == 32'h02000040));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004008) == 32'h00004008));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL_1 = (|{((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002040) == 32'h00002040),((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001040) == 32'h00001040)});
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004000) == 32'h00004000));
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK_2 = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_2 = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1 = 1'b0;
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO_1 = (|((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000008) == 32'h00000008));
  assign _zz_DispatchPlugin_logic_ptr_next = (CommitPlugin_logic_commit_reschedulePort_payload_robIdNext - 6'h20);
  assign _zz_DispatchPlugin_logic_push_commitNotWaitingOnUs = ((CommitPlugin_logic_commit_head ^ FrontendPlugin_dispatch_ROB_ID) >>> 1'd1);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_0 = (32'h00000001 <<< _zz_DispatchPlugin_logic_push_slots_0_events_0_1);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_0_2 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0 - DispatchPlugin_logic_ptr_next);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_0_1 = _zz_DispatchPlugin_logic_push_slots_0_events_0_2[4:0];
  assign _zz_DispatchPlugin_logic_push_slots_0_events_1 = (32'h00000001 <<< _zz_DispatchPlugin_logic_push_slots_0_events_1_1);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_1_2 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0 - DispatchPlugin_logic_ptr_next);
  assign _zz_DispatchPlugin_logic_push_slots_0_events_1_1 = _zz_DispatchPlugin_logic_push_slots_0_events_1_2[4:0];
  assign _zz_DispatchPlugin_logic_push_slots_1_events_0 = (32'h00000001 <<< _zz_DispatchPlugin_logic_push_slots_1_events_0_1);
  assign _zz_DispatchPlugin_logic_push_slots_1_events_0_2 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_1 - DispatchPlugin_logic_ptr_next);
  assign _zz_DispatchPlugin_logic_push_slots_1_events_0_1 = _zz_DispatchPlugin_logic_push_slots_1_events_0_2[4:0];
  assign _zz_DispatchPlugin_logic_push_slots_1_events_1 = (32'h00000001 <<< _zz_DispatchPlugin_logic_push_slots_1_events_1_1);
  assign _zz_DispatchPlugin_logic_push_slots_1_events_1_2 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_1 - DispatchPlugin_logic_ptr_next);
  assign _zz_DispatchPlugin_logic_push_slots_1_events_1_1 = _zz_DispatchPlugin_logic_push_slots_1_events_1_2[4:0];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID = {1'd0, DispatchPlugin_logic_pop_0_stagesList_1_UINT};
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID = {1'd0, DispatchPlugin_logic_pop_1_stagesList_1_UINT};
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_1_ROB_ID = {1'd0, DispatchPlugin_logic_pop_2_stagesList_1_UINT};
  assign _zz_DispatchPlugin_logic_wake_dynamic_offseted_0_payload = (Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_payload_robId - DispatchPlugin_logic_ptr_current);
  assign _zz_DispatchPlugin_logic_wake_dynamic_offseted_1_payload = (Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_payload_robId - DispatchPlugin_logic_ptr_current);
  assign _zz_DispatchPlugin_logic_wake_dynamic_offseted_2_payload = (Lsu2Plugin_logic_special_wakeRob_payload_robId - DispatchPlugin_logic_ptr_current);
  assign _zz_DispatchPlugin_logic_wake_dynamic_offseted_3_payload = (EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_payload_robId - DispatchPlugin_logic_ptr_current);
  assign _zz_DispatchPlugin_logic_wake_dynamic_masks_0 = (32'h00000001 <<< DispatchPlugin_logic_wake_dynamic_offseted_0_payload);
  assign _zz_DispatchPlugin_logic_wake_dynamic_masks_1 = (32'h00000001 <<< DispatchPlugin_logic_wake_dynamic_offseted_1_payload);
  assign _zz_DispatchPlugin_logic_wake_dynamic_masks_2 = (32'h00000001 <<< DispatchPlugin_logic_wake_dynamic_offseted_2_payload);
  assign _zz_DispatchPlugin_logic_wake_dynamic_masks_3 = (32'h00000001 <<< DispatchPlugin_logic_wake_dynamic_offseted_3_payload);
  assign _zz_RobPlugin_logic_completionMem_init_0_robId = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_RobPlugin_logic_completionMem_init_1_robId = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz__zz_CommitPlugin_setup_robLineMask_mask = (CommitPlugin_setup_robLineMask_line >>> 1'd1);
  assign _zz__zz_CommitPlugin_setup_robLineMask_mask_1 = (CommitPlugin_setup_robLineMask_line >>> 1'd1);
  assign _zz__zz_when_RobPlugin_l118 = (CommitPlugin_setup_robLineMask_line >>> 1'd1);
  assign _zz__zz_when_RobPlugin_l118_1 = (CommitPlugin_setup_robLineMask_line >>> 1'd1);
  assign _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz__zz_CommitPlugin_logic_commit_active_2 = {_zz_CommitPlugin_logic_commit_active_1[1],_zz_CommitPlugin_logic_commit_active_1[0]};
  assign _zz__zz_integer_RfAllocationPlugin_logic_push_mask_0_2 = {_zz_integer_RfAllocationPlugin_logic_push_mask_0_1[1],_zz_integer_RfAllocationPlugin_logic_push_mask_0_1[0]};
  assign _zz__zz_commit_pc_0_1 = {_zz_RobPlugin_logic_storage_PC_banks_1_port1[31 : 0],_zz_RobPlugin_logic_storage_PC_banks_0_port1[31 : 0]};
  assign _zz__zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1 = {_zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port1[0],_zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port1[0]};
  assign _zz__zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1 = {_zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port2[0],_zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port2[0]};
  assign _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz__zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2 = {_zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_1[11 : 6],_zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_1[5 : 0]};
  assign _zz__zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2 = {_zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_1[11 : 6],_zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_1[5 : 0]};
  assign _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz__zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2 = {_zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_1[9 : 5],_zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_1[4 : 0]};
  assign _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz__zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2 = {_zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_1[11 : 6],_zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_1[5 : 0]};
  assign _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz__zz_BranchContextPlugin_logic_onCommit_isBranch_0_2 = {_zz_BranchContextPlugin_logic_onCommit_isBranch_0_1[1],_zz_BranchContextPlugin_logic_onCommit_isBranch_0_1[0]};
  assign _zz__zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1 = {_zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port1[0],_zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port1[0]};
  assign _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port = (FrontendPlugin_dispatch_ROB_ID >>> 1'd1);
  assign _zz__zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2 = {_zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_1[1],_zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_1[0]};
  assign _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port = (FrontendPlugin_dispatch_ROB_ID >>> 1'd1);
  assign _zz__zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2 = {_zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_1[1],_zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_1[0]};
  assign _zz_PcPlugin_logic_init_counter_1 = (! PcPlugin_logic_init_booted);
  assign _zz_PcPlugin_logic_init_counter = {6'd0, _zz_PcPlugin_logic_init_counter_1};
  assign _zz_PcPlugin_logic_fetchPc_pc_1 = ({3'd0,PcPlugin_logic_fetchPc_inc} <<< 2'd3);
  assign _zz_PcPlugin_logic_fetchPc_pc = {28'd0, _zz_PcPlugin_logic_fetchPc_pc_1};
  assign _zz_PerformanceCounterPlugin_setup_writePort_data = PerformanceCounterPlugin_logic_fsm_result;
  assign _zz_PerformanceCounterPlugin_setup_writePort_data_1 = (PerformanceCounterPlugin_logic_fsm_result >>> 6'd32);
  assign _zz_PerformanceCounterPlugin_setup_writePort_address_1 = {2'd0, PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address};
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2_1 = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3_2 = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4_2 = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5_2 = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6_2 = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign _zz_PrivilegedPlugin_setup_ramWrite_data = PrivilegedPlugin_logic_reschedule_payload_epc;
  assign _zz_PrivilegedPlugin_setup_ramWrite_data_1 = PrivilegedPlugin_logic_reschedule_payload_tval;
  assign _zz_PrivilegedPlugin_logic_readed = (PrivilegedPlugin_logic_reschedule_payload_epc + _zz_PrivilegedPlugin_logic_readed_1);
  assign _zz_PrivilegedPlugin_logic_readed_2 = ((PrivilegedPlugin_logic_reschedule_payload_cause != 4'b1010) ? _zz_PrivilegedPlugin_logic_readed_3 : 4'b0000);
  assign _zz_PrivilegedPlugin_logic_readed_1 = {28'd0, _zz_PrivilegedPlugin_logic_readed_2};
  assign _zz_PrivilegedPlugin_logic_readed_3 = ({2'd0,_zz_PrivilegedPlugin_logic_readed_4} <<< 2'd2);
  assign _zz_PrivilegedPlugin_logic_readed_4 = (_zz_PrivilegedPlugin_logic_readed_5 + {1'b0,1'b1});
  assign _zz_PrivilegedPlugin_logic_readed_6 = 1'b0;
  assign _zz_PrivilegedPlugin_logic_readed_5 = {1'd0, _zz_PrivilegedPlugin_logic_readed_6};
  assign _zz_FetchCachePlugin_logic_ways_0_mem_port = {FetchCachePlugin_logic_waysWrite_tag_address,{FetchCachePlugin_logic_waysWrite_tag_error,FetchCachePlugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchCachePlugin_logic_ways_0_mem_port_1 = FetchCachePlugin_logic_waysWrite_mask[0];
  assign _zz_FetchCachePlugin_logic_ways_1_mem_port = {FetchCachePlugin_logic_waysWrite_tag_address,{FetchCachePlugin_logic_waysWrite_tag_error,FetchCachePlugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchCachePlugin_logic_ways_1_mem_port_1 = FetchCachePlugin_logic_waysWrite_mask[1];
  assign _zz_FetchCachePlugin_logic_ways_2_mem_port = {FetchCachePlugin_logic_waysWrite_tag_address,{FetchCachePlugin_logic_waysWrite_tag_error,FetchCachePlugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchCachePlugin_logic_ways_2_mem_port_1 = FetchCachePlugin_logic_waysWrite_mask[2];
  assign _zz_FetchCachePlugin_logic_ways_3_mem_port = {FetchCachePlugin_logic_waysWrite_tag_address,{FetchCachePlugin_logic_waysWrite_tag_error,FetchCachePlugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchCachePlugin_logic_ways_3_mem_port_1 = FetchCachePlugin_logic_waysWrite_mask[3];
  assign _zz_FetchCachePlugin_logic_plru_ram_port = {FetchCachePlugin_logic_plru_write_payload_data_1,FetchCachePlugin_logic_plru_write_payload_data_0};
  assign _zz_DecoderPredictionPlugin_logic_ras_mem_stack_port = DecoderPredictionPlugin_logic_ras_write_payload_data;
  assign _zz_BtbPlugin_logic_mem_port = {BtbPlugin_logic_onLearn_port_payload_data_isBranch,{BtbPlugin_logic_onLearn_port_payload_data_pcTarget,{BtbPlugin_logic_onLearn_port_payload_data_slice,BtbPlugin_logic_onLearn_port_payload_data_hash}}};
  assign _zz_GSharePlugin_logic_mem_counter_port = {GSharePlugin_logic_mem_write_payload_data_1,GSharePlugin_logic_mem_write_payload_data_0};
  assign _zz_Lsu2Plugin_logic_lq_mem_addressPre_port_1 = AguPlugin_setup_port_payload_address;
  assign _zz_Lsu2Plugin_logic_lq_mem_addressPost_port = Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
  assign _zz_Lsu2Plugin_logic_lq_mem_size_port_1 = AguPlugin_setup_port_payload_size;
  assign _zz_Lsu2Plugin_logic_lq_mem_physRd_port_1 = AguPlugin_setup_port_payload_physicalRd;
  assign _zz_Lsu2Plugin_logic_lq_mem_robId_port_1 = AguPlugin_setup_port_payload_robId;
  assign _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port_1 = AguPlugin_setup_port_payload_robIdMsb;
  assign _zz_Lsu2Plugin_logic_lq_mem_pc_port_1 = AguPlugin_setup_port_payload_pc;
  assign _zz_Lsu2Plugin_logic_lq_mem_io_port = Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO;
  assign _zz_Lsu2Plugin_logic_lq_mem_writeRd_port_1 = AguPlugin_setup_port_payload_writeRd;
  assign _zz_Lsu2Plugin_logic_lq_mem_lr_port_1 = AguPlugin_setup_port_payload_lr;
  assign _zz_Lsu2Plugin_logic_lq_mem_unsigned_port_1 = AguPlugin_setup_port_payload_unsigned;
  assign _zz_Lsu2Plugin_logic_lq_mem_spFpAddress_port = ({(FrontendPlugin_dispatch_ARCH_RS_0_0 == 5'h08),{(FrontendPlugin_dispatch_ARCH_RS_0_0 == 5'h03),(FrontendPlugin_dispatch_ARCH_RS_0_0 == 5'h02)}} != 3'b000);
  assign _zz_Lsu2Plugin_logic_lq_mem_spFpAddress_port_1 = ({(FrontendPlugin_dispatch_ARCH_RS_0_1 == 5'h08),{(FrontendPlugin_dispatch_ARCH_RS_0_1 == 5'h03),(FrontendPlugin_dispatch_ARCH_RS_0_1 == 5'h02)}} != 3'b000);
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port_1 = Lsu2Plugin_logic_aguPush_0_hazardPrediction_hit;
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port_1 = Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_delta;
  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port_1 = Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
  assign _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port_1 = Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter;
  assign _zz_Lsu2Plugin_logic_sq_mem_robId_port_1 = AguPlugin_setup_port_payload_robId;
  assign _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port_1 = AguPlugin_setup_port_payload_robIdMsb;
  assign _zz_Lsu2Plugin_logic_sq_mem_addressPre_port_1 = AguPlugin_setup_port_payload_address;
  assign _zz_Lsu2Plugin_logic_sq_mem_addressPost_port = Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
  assign _zz_Lsu2Plugin_logic_sq_mem_size_port_1 = AguPlugin_setup_port_payload_size;
  assign _zz_Lsu2Plugin_logic_sq_mem_io_port = Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO;
  assign _zz_Lsu2Plugin_logic_sq_mem_amo_port_1 = AguPlugin_setup_port_payload_amo;
  assign _zz_Lsu2Plugin_logic_sq_mem_sc_port_1 = AguPlugin_setup_port_payload_sc;
  assign _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port_1 = (AguPlugin_setup_port_payload_amo || AguPlugin_setup_port_payload_sc);
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port = {FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask[0];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port = {FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask[1];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port = {FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask[2];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port = {FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask[3];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port = {FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask[0];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port = {FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault,{FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault,FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid}}}}}}}};
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port_1 = FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask[1];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port = {Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask[0];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port = {Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask[1];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port = {Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask[2];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port = {Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask[3];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port = {Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask[0];
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port = {Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault,{Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault,Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid}}}}}}}};
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port_1 = Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask[1];
  assign _zz_RobPlugin_logic_completionMem_hits_0_port = (! _zz_RobPlugin_logic_completionMem_hits_0_port2[0]);
  assign _zz_RobPlugin_logic_completionMem_hits_1_port = (! _zz_RobPlugin_logic_completionMem_hits_1_port2[0]);
  assign _zz_RobPlugin_logic_completionMem_hits_2_port = (! _zz_RobPlugin_logic_completionMem_hits_2_port2[0]);
  assign _zz_RobPlugin_logic_completionMem_hits_3_port = (! _zz_RobPlugin_logic_completionMem_hits_3_port2[0]);
  assign _zz_RobPlugin_logic_completionMem_hits_4_port = (! _zz_RobPlugin_logic_completionMem_hits_4_port2[0]);
  assign _zz_RobPlugin_logic_completionMem_hits_5_port = (! _zz_RobPlugin_logic_completionMem_hits_5_port2[0]);
  assign _zz_RobPlugin_logic_completionMem_hits_6_port = (! _zz_RobPlugin_logic_completionMem_hits_6_port2[0]);
  assign _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port_1 = {FrontendPlugin_allocated_Frontend_DISPATCH_MASK_1,FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0};
  assign _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port_2 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PC_banks_0_port = FrontendPlugin_allocated_PC_0;
  assign _zz_RobPlugin_logic_storage_PC_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PC_banks_1_port = FrontendPlugin_allocated_PC_1;
  assign _zz_RobPlugin_logic_storage_PC_banks_1_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port = FrontendPlugin_allocated_WRITE_RD_0;
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port = FrontendPlugin_allocated_WRITE_RD_1;
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port_1 = {FrontendPlugin_allocated_PHYS_RD_1,FrontendPlugin_allocated_PHYS_RD_0};
  assign _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port_2 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port_1 = {FrontendPlugin_allocated_ARCH_RD_1,FrontendPlugin_allocated_ARCH_RD_0};
  assign _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port_2 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port_1 = {FrontendPlugin_allocated_PHYS_RD_FREE_1,FrontendPlugin_allocated_PHYS_RD_FREE_0};
  assign _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port_2 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port_1 = {FrontendPlugin_allocated_BRANCH_SEL_1,FrontendPlugin_allocated_BRANCH_SEL_0};
  assign _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port_2 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port = FrontendPlugin_dispatch_Prediction_IS_BRANCH_0;
  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port_1 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port = FrontendPlugin_dispatch_Prediction_IS_BRANCH_1;
  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port_1 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_port = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_1_port = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port = FrontendPlugin_allocated_DecoderPredictionPlugin_RAS_PUSH_PTR_0;
  assign _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1_port = FrontendPlugin_allocated_DecoderPredictionPlugin_RAS_PUSH_PTR_1;
  assign _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port_1 = {FrontendPlugin_dispatch_LQ_ALLOC_1,FrontendPlugin_dispatch_LQ_ALLOC_0};
  assign _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port_2 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port_1 = {FrontendPlugin_dispatch_SQ_ALLOC_1,FrontendPlugin_dispatch_SQ_ALLOC_0};
  assign _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port_2 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1_port = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port = FrontendPlugin_allocated_PHYS_RS_0_0;
  assign _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_1_port = FrontendPlugin_allocated_PHYS_RS_0_1;
  assign _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_1_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port = FrontendPlugin_allocated_READ_RS_0_0;
  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port = FrontendPlugin_allocated_READ_RS_0_1;
  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port = FrontendPlugin_allocated_PHYS_RS_1_0;
  assign _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_1_port = FrontendPlugin_allocated_PHYS_RS_1_1;
  assign _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_1_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port = FrontendPlugin_allocated_READ_RS_1_0;
  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port = FrontendPlugin_allocated_READ_RS_1_1;
  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port = FrontendPlugin_allocated_BRANCH_ID_0;
  assign _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_BRANCH_ID_banks_1_port = FrontendPlugin_allocated_BRANCH_ID_1;
  assign _zz_RobPlugin_logic_storage_BRANCH_ID_banks_1_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port = FrontendPlugin_dispatch_LSU_ID_0;
  assign _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port_1 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_LSU_ID_banks_1_port = FrontendPlugin_dispatch_LSU_ID_1;
  assign _zz_RobPlugin_logic_storage_LSU_ID_banks_1_port_1 = (FrontendPlugin_dispatch_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port = FrontendPlugin_allocated_ROB_MSB_0;
  assign _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_RobPlugin_logic_storage_ROB_MSB_banks_1_port = FrontendPlugin_allocated_ROB_MSB_1;
  assign _zz_RobPlugin_logic_storage_ROB_MSB_banks_1_port_1 = (FrontendPlugin_allocated_isFireing && 1'b1);
  assign _zz_FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT_1 = FetchPlugin_stages_1_Fetch_FETCH_PC[2 : 2];
  assign _zz_AlignerPlugin_logic_extractors_0_pcWord_1 = AlignerPlugin_logic_extractors_0_firstWord;
  assign _zz_AlignerPlugin_logic_extractors_1_pcWord_1 = AlignerPlugin_logic_extractors_1_firstWord;
  assign _zz_CommitDebugFilterPlugin_logic_commits_3 = {_zz_CommitDebugFilterPlugin_logic_commits_1,_zz_CommitDebugFilterPlugin_logic_commits};
  assign _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_3 = CommitPlugin_logic_commit_reschedulePort_payload_robId[0 : 0];
  assign _zz_PerformanceCounterPlugin_logic_commitCount_1 = {_zz_CommitDebugFilterPlugin_logic_commits_1,_zz_CommitDebugFilterPlugin_logic_commits};
  assign _zz_PerformanceCounterPlugin_logic_events_sums_0_1 = FetchCachePlugin_setup_refillEvent;
  assign _zz_PerformanceCounterPlugin_logic_events_sums_1_1 = DataCachePlugin_setup_refillEvent;
  assign _zz_PerformanceCounterPlugin_logic_events_sums_2_1 = DataCachePlugin_setup_writebackEvent;
  assign _zz_PerformanceCounterPlugin_logic_events_sums_3_1 = PerformanceCounterPlugin_logic_branchMissEvent;
  assign _zz_BranchContextPlugin_logic_onCommit_commitedNext_2 = {BranchContextPlugin_logic_onCommit_isBranchCommit_1,BranchContextPlugin_logic_onCommit_isBranchCommit_0};
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_3 = CommitPlugin_logic_reschedule_reschedulePort_payload_robId[0 : 0];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_3 = CommitPlugin_logic_reschedule_reschedulePort_payload_robId[0 : 0];
  assign _zz_DecoderPredictionPlugin_logic_ras_healPush_3 = CommitPlugin_logic_reschedule_reschedulePort_payload_robId[0 : 0];
  assign _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount_1 = {Lsu2Plugin_logic_lq_onCommit_lqCommits_1,Lsu2Plugin_logic_lq_onCommit_lqCommits_0};
  assign _zz_Lsu2Plugin_logic_allocation_loads_requestsCount_1 = {Lsu2Plugin_logic_allocation_loads_requests_1,Lsu2Plugin_logic_allocation_loads_requests_0};
  assign _zz_Lsu2Plugin_logic_allocation_stores_requestsCount_1 = {Lsu2Plugin_logic_allocation_stores_requests_1,Lsu2Plugin_logic_allocation_stores_requests_0};
  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_1 = Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress[1 : 0];
  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_3 = Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress[1 : 1];
  assign _zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17_1 = EU0_CsrAccessPlugin_setup_onReadAddress[7];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_3 = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_3 = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_3 = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_3 = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_3 = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_3 = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID[0 : 0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_3 = EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID[0 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_3 = {_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1,_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data};
  assign _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_3 = {_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1,_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data};
  assign _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_3 = {_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1,_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data};
  assign _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_3 = {_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1,_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data};
  assign _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_3 = {_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1,_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data};
  assign _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_3 = {_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1,_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data};
  assign _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_1 = _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[6];
  assign _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_2 = _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[7];
  assign _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_3 = {_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[8],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[9],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[10],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[11],_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[12]}}}};
  assign _zz_GSharePlugin_logic_onLearn_hash_1 = _zz_GSharePlugin_logic_onLearn_hash[6];
  assign _zz_GSharePlugin_logic_onLearn_hash_2 = _zz_GSharePlugin_logic_onLearn_hash[7];
  assign _zz_GSharePlugin_logic_onLearn_hash_3 = {_zz_GSharePlugin_logic_onLearn_hash[8],{_zz_GSharePlugin_logic_onLearn_hash[9],{_zz_GSharePlugin_logic_onLearn_hash[10],{_zz_GSharePlugin_logic_onLearn_hash[11],_zz_GSharePlugin_logic_onLearn_hash[12]}}}};
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits = (! CommitPlugin_logic_reschedule_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_1 = (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age < CommitPlugin_logic_reschedule_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_2 = (! Lsu2Plugin_setup_specialTrap_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_3 = (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_1_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_4 = (! CommitPlugin_logic_reschedule_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_5 = (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age < CommitPlugin_logic_reschedule_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_6 = (! Lsu2Plugin_setup_sharedTrap_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_7 = (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age < CommitPlugin_logic_reschedule_portsLogic_perPort_0_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_8 = (! CommitPlugin_logic_reschedule_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_9 = (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age < CommitPlugin_logic_reschedule_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_10 = (! Lsu2Plugin_setup_sharedTrap_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_11 = (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age < CommitPlugin_logic_reschedule_portsLogic_perPort_0_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_12 = (! CommitPlugin_logic_reschedule_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_13 = (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_age);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_14 = (! Lsu2Plugin_setup_sharedTrap_valid);
  assign _zz_CommitPlugin_logic_reschedule_portsLogic_hits_15 = (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_portsLogic_perPort_0_age);
  assign _zz_CommitPlugin_logic_reschedule_robId = Lsu2Plugin_setup_sharedTrap_payload_robId;
  assign _zz_CommitPlugin_logic_reschedule_robId_1 = 6'h00;
  assign _zz_CommitPlugin_logic_reschedule_robId_2 = Lsu2Plugin_setup_specialTrap_payload_robId;
  assign _zz_CommitPlugin_logic_reschedule_robId_3 = 6'h00;
  assign _zz_CommitPlugin_logic_reschedule_robId_4 = ALU0_BranchPlugin_setup_reschedule_payload_robId;
  assign _zz_CommitPlugin_logic_reschedule_robId_5 = 6'h00;
  assign _zz_CommitPlugin_logic_reschedule_robId_6 = EnvCallPlugin_setup_reschedule_payload_robId;
  assign _zz_CommitPlugin_logic_reschedule_robId_7 = 6'h00;
  assign _zz_CommitPlugin_logic_reschedule_cause = CommitPlugin_logic_reschedule_portsLogic_hits[0];
  assign _zz_CommitPlugin_logic_reschedule_cause_1 = Lsu2Plugin_setup_sharedTrap_payload_cause;
  assign _zz_CommitPlugin_logic_reschedule_cause_2 = 4'b0000;
  assign _zz_CommitPlugin_logic_reschedule_cause_3 = CommitPlugin_logic_reschedule_portsLogic_hits[1];
  assign _zz_CommitPlugin_logic_reschedule_cause_4 = Lsu2Plugin_setup_specialTrap_payload_cause;
  assign _zz_CommitPlugin_logic_reschedule_cause_5 = 4'b0000;
  assign _zz_CommitPlugin_logic_reschedule_cause_6 = CommitPlugin_logic_reschedule_portsLogic_hits[2];
  assign _zz_CommitPlugin_logic_reschedule_cause_7 = ALU0_BranchPlugin_setup_reschedule_payload_cause;
  assign _zz_CommitPlugin_logic_reschedule_cause_8 = 4'b0000;
  assign _zz_CommitPlugin_logic_reschedule_cause_9 = CommitPlugin_logic_reschedule_portsLogic_hits[3];
  assign _zz_CommitPlugin_logic_reschedule_cause_10 = EnvCallPlugin_setup_reschedule_payload_cause;
  assign _zz_CommitPlugin_logic_reschedule_cause_11 = 4'b0000;
  assign _zz_CommitPlugin_logic_reschedule_reason = CommitPlugin_logic_reschedule_portsLogic_hits[0];
  assign _zz_CommitPlugin_logic_reschedule_reason_1 = Lsu2Plugin_setup_sharedTrap_payload_reason;
  assign _zz_CommitPlugin_logic_reschedule_reason_2 = 8'h00;
  assign _zz_CommitPlugin_logic_reschedule_reason_3 = CommitPlugin_logic_reschedule_portsLogic_hits[1];
  assign _zz_CommitPlugin_logic_reschedule_reason_4 = Lsu2Plugin_setup_specialTrap_payload_reason;
  assign _zz_CommitPlugin_logic_reschedule_reason_5 = 8'h00;
  assign _zz_CommitPlugin_logic_reschedule_reason_6 = CommitPlugin_logic_reschedule_portsLogic_hits[2];
  assign _zz_CommitPlugin_logic_reschedule_reason_7 = ALU0_BranchPlugin_setup_reschedule_payload_reason;
  assign _zz_CommitPlugin_logic_reschedule_reason_8 = 8'h00;
  assign _zz_CommitPlugin_logic_reschedule_reason_9 = CommitPlugin_logic_reschedule_portsLogic_hits[3];
  assign _zz_CommitPlugin_logic_reschedule_reason_10 = EnvCallPlugin_setup_reschedule_payload_reason;
  assign _zz_CommitPlugin_logic_reschedule_reason_11 = 8'h00;
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_1 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[9];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_2 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[10];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_3 = {ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[11],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[12],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[13],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[14],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[15],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[16],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[17],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[18],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[19],{_zz_ALU0_ShiftPlugin_logic_process_reversed_4,{_zz_ALU0_ShiftPlugin_logic_process_reversed_5,_zz_ALU0_ShiftPlugin_logic_process_reversed_6}}}}}}}}}}};
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_4 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[20];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_5 = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[21];
  assign _zz_ALU0_ShiftPlugin_logic_process_reversed_6 = {ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[22],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[23],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[24],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[25],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[26],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[27],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[28],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[29],{ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[30],ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]}}}}}}}}};
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_1 = ALU0_ShiftPlugin_logic_process_shifted[9];
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_2 = ALU0_ShiftPlugin_logic_process_shifted[10];
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_3 = {ALU0_ShiftPlugin_logic_process_shifted[11],{ALU0_ShiftPlugin_logic_process_shifted[12],{ALU0_ShiftPlugin_logic_process_shifted[13],{ALU0_ShiftPlugin_logic_process_shifted[14],{ALU0_ShiftPlugin_logic_process_shifted[15],{ALU0_ShiftPlugin_logic_process_shifted[16],{ALU0_ShiftPlugin_logic_process_shifted[17],{ALU0_ShiftPlugin_logic_process_shifted[18],{ALU0_ShiftPlugin_logic_process_shifted[19],{_zz_ALU0_ShiftPlugin_logic_process_patched_4,{_zz_ALU0_ShiftPlugin_logic_process_patched_5,_zz_ALU0_ShiftPlugin_logic_process_patched_6}}}}}}}}}}};
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_4 = ALU0_ShiftPlugin_logic_process_shifted[20];
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_5 = ALU0_ShiftPlugin_logic_process_shifted[21];
  assign _zz_ALU0_ShiftPlugin_logic_process_patched_6 = {ALU0_ShiftPlugin_logic_process_shifted[22],{ALU0_ShiftPlugin_logic_process_shifted[23],{ALU0_ShiftPlugin_logic_process_shifted[24],{ALU0_ShiftPlugin_logic_process_shifted[25],{ALU0_ShiftPlugin_logic_process_shifted[26],{ALU0_ShiftPlugin_logic_process_shifted[27],{ALU0_ShiftPlugin_logic_process_shifted[28],{ALU0_ShiftPlugin_logic_process_shifted[29],{ALU0_ShiftPlugin_logic_process_shifted[30],ALU0_ShiftPlugin_logic_process_shifted[31]}}}}}}}}};
  assign _zz_ALU1_ShiftPlugin_logic_process_reversed_1 = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[9];
  assign _zz_ALU1_ShiftPlugin_logic_process_reversed_2 = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[10];
  assign _zz_ALU1_ShiftPlugin_logic_process_reversed_3 = {ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[11],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[12],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[13],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[14],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[15],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[16],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[17],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[18],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[19],{_zz_ALU1_ShiftPlugin_logic_process_reversed_4,{_zz_ALU1_ShiftPlugin_logic_process_reversed_5,_zz_ALU1_ShiftPlugin_logic_process_reversed_6}}}}}}}}}}};
  assign _zz_ALU1_ShiftPlugin_logic_process_reversed_4 = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[20];
  assign _zz_ALU1_ShiftPlugin_logic_process_reversed_5 = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[21];
  assign _zz_ALU1_ShiftPlugin_logic_process_reversed_6 = {ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[22],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[23],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[24],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[25],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[26],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[27],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[28],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[29],{ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[30],ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]}}}}}}}}};
  assign _zz_ALU1_ShiftPlugin_logic_process_patched_1 = ALU1_ShiftPlugin_logic_process_shifted[9];
  assign _zz_ALU1_ShiftPlugin_logic_process_patched_2 = ALU1_ShiftPlugin_logic_process_shifted[10];
  assign _zz_ALU1_ShiftPlugin_logic_process_patched_3 = {ALU1_ShiftPlugin_logic_process_shifted[11],{ALU1_ShiftPlugin_logic_process_shifted[12],{ALU1_ShiftPlugin_logic_process_shifted[13],{ALU1_ShiftPlugin_logic_process_shifted[14],{ALU1_ShiftPlugin_logic_process_shifted[15],{ALU1_ShiftPlugin_logic_process_shifted[16],{ALU1_ShiftPlugin_logic_process_shifted[17],{ALU1_ShiftPlugin_logic_process_shifted[18],{ALU1_ShiftPlugin_logic_process_shifted[19],{_zz_ALU1_ShiftPlugin_logic_process_patched_4,{_zz_ALU1_ShiftPlugin_logic_process_patched_5,_zz_ALU1_ShiftPlugin_logic_process_patched_6}}}}}}}}}}};
  assign _zz_ALU1_ShiftPlugin_logic_process_patched_4 = ALU1_ShiftPlugin_logic_process_shifted[20];
  assign _zz_ALU1_ShiftPlugin_logic_process_patched_5 = ALU1_ShiftPlugin_logic_process_shifted[21];
  assign _zz_ALU1_ShiftPlugin_logic_process_patched_6 = {ALU1_ShiftPlugin_logic_process_shifted[22],{ALU1_ShiftPlugin_logic_process_shifted[23],{ALU1_ShiftPlugin_logic_process_shifted[24],{ALU1_ShiftPlugin_logic_process_shifted[25],{ALU1_ShiftPlugin_logic_process_shifted[26],{ALU1_ShiftPlugin_logic_process_shifted[27],{ALU1_ShiftPlugin_logic_process_shifted[28],{ALU1_ShiftPlugin_logic_process_shifted[29],{ALU1_ShiftPlugin_logic_process_shifted[30],ALU1_ShiftPlugin_logic_process_shifted[31]}}}}}}}}};
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo = Lsu2Plugin_logic_lq_regs_5_redo;
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_1 = {Lsu2Plugin_logic_lq_regs_4_redo,{Lsu2Plugin_logic_lq_regs_3_redo,{Lsu2Plugin_logic_lq_regs_2_redo,{Lsu2Plugin_logic_lq_regs_1_redo,Lsu2Plugin_logic_lq_regs_0_redo}}}};
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo = Lsu2Plugin_logic_sq_regs_5_redo;
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_1 = {Lsu2Plugin_logic_sq_regs_4_redo,{Lsu2Plugin_logic_sq_regs_3_redo,{Lsu2Plugin_logic_sq_regs_2_redo,{Lsu2Plugin_logic_sq_regs_1_redo,Lsu2Plugin_logic_sq_regs_0_redo}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_1 = 4'b1010;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_2 = (4'b1001 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_3 = (4'b1000 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_4 = {(4'b0111 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(4'b0110 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(4'b0101 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(4'b0100 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(4'b0011 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(4'b0010 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_5 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),(_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_6 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask)}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_5 = 4'b0001;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_6 = 4'b0000;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_1 = 4'b1010;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_2 = (4'b1001 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_3 = (4'b1000 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_4 = {(4'b0111 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(4'b0110 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(4'b0101 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(4'b0100 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(4'b0011 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(4'b0010 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_5 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),(_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_6 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask)}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_5 = 4'b0001;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_6 = 4'b0000;
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input_1 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[7];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input_2 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[8];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input_3 = {_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[9],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[10],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[11],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[12],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[13],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[14],_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[15]}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits_1 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[7];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits_2 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[8];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits_3 = {_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[9],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[10],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[11],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[12],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[13],_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[14]}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[7];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh_1 = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[8];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh_2 = {Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[9],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[10],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[11],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[12],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[13],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[14],Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[15]}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_1 = 4'b1010;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_2 = (4'b1001 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_3 = (4'b1000 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_4 = {(4'b0111 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(4'b0110 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(4'b0101 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(4'b0100 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(4'b0011 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(4'b0010 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_5 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),(_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_6 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask)}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_5 = 4'b0001;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_6 = 4'b0000;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_1 = 4'b1010;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_2 = (4'b1001 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_3 = (4'b1000 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_4 = {(4'b0111 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(4'b0110 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(4'b0101 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(4'b0100 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(4'b0011 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(4'b0010 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_5 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),(_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_6 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask)}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_5 = 4'b0001;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_6 = 4'b0000;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_physicalAddress,_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_1};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_2 = 32'h00000000;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_3 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_physicalAddress,_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_4};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_5 = 32'h00000000;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_6 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_physicalAddress,_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_7};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_8 = 32'h00000000;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_9 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_physicalAddress,_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_10};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_11 = 32'h00000000;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_12 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[21 : 0]};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_13 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[21 : 0]};
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_1 = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_4 = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_7 = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_10 = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated = {FetchPlugin_stages_1_MMU_L0_ENTRIES_0_physicalAddress,_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_1};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_2 = 32'h00000000;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_3 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_1_physicalAddress,_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_4};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_5 = 32'h00000000;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_6 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_2_physicalAddress,_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_7};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_8 = 32'h00000000;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_9 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_3_physicalAddress,_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_10};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_11 = 32'h00000000;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_12 = {FetchPlugin_stages_1_MMU_L1_ENTRIES_0_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[21 : 0]};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_13 = {FetchPlugin_stages_1_MMU_L1_ENTRIES_1_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[21 : 0]};
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_1 = FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_4 = FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_7 = FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_10 = FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0];
  assign _zz_COMB_CSR_ = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__1 = 12'hb9e;
  assign _zz_COMB_CSR__2 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb1e);
  assign _zz_COMB_CSR__3 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h33d);
  assign _zz_COMB_CSR__4 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb9d),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb1d),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h33c),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb9c),{(_zz_COMB_CSR__5 == _zz_COMB_CSR__6),{_zz_COMB_CSR__7,{_zz_COMB_CSR__8,_zz_COMB_CSR__9}}}}}}};
  assign _zz_COMB_CSR__5 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__6 = 12'hb1c;
  assign _zz_COMB_CSR__7 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h33b);
  assign _zz_COMB_CSR__8 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb9b);
  assign _zz_COMB_CSR__9 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb1b),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h33a),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb9a),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb1a),{(_zz_COMB_CSR__10 == _zz_COMB_CSR__11),{_zz_COMB_CSR__12,{_zz_COMB_CSR__13,_zz_COMB_CSR__14}}}}}}};
  assign _zz_COMB_CSR__10 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__11 = 12'h339;
  assign _zz_COMB_CSR__12 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb99);
  assign _zz_COMB_CSR__13 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb19);
  assign _zz_COMB_CSR__14 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h338),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb98),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb18),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h337),{(_zz_COMB_CSR__15 == _zz_COMB_CSR__16),{_zz_COMB_CSR__17,{_zz_COMB_CSR__18,_zz_COMB_CSR__19}}}}}}};
  assign _zz_COMB_CSR__15 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__16 = 12'hb97;
  assign _zz_COMB_CSR__17 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb17);
  assign _zz_COMB_CSR__18 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h336);
  assign _zz_COMB_CSR__19 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb96),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb16),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h335),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb95),{(_zz_COMB_CSR__20 == _zz_COMB_CSR__21),{_zz_COMB_CSR__22,{_zz_COMB_CSR__23,_zz_COMB_CSR__24}}}}}}};
  assign _zz_COMB_CSR__20 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__21 = 12'hb15;
  assign _zz_COMB_CSR__22 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h334);
  assign _zz_COMB_CSR__23 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb94);
  assign _zz_COMB_CSR__24 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb14),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h333),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb93),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb13),{(_zz_COMB_CSR__25 == _zz_COMB_CSR__26),{_zz_COMB_CSR__27,{_zz_COMB_CSR__28,_zz_COMB_CSR__29}}}}}}};
  assign _zz_COMB_CSR__25 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__26 = 12'h332;
  assign _zz_COMB_CSR__27 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb92);
  assign _zz_COMB_CSR__28 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb12);
  assign _zz_COMB_CSR__29 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h331),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb91),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb11),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h330),{(_zz_COMB_CSR__30 == _zz_COMB_CSR__31),{_zz_COMB_CSR__32,{_zz_COMB_CSR__33,_zz_COMB_CSR__34}}}}}}};
  assign _zz_COMB_CSR__30 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__31 = 12'hb90;
  assign _zz_COMB_CSR__32 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb10);
  assign _zz_COMB_CSR__33 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h32f);
  assign _zz_COMB_CSR__34 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb8f),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb0f),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h32e),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb8e),{(_zz_COMB_CSR__35 == _zz_COMB_CSR__36),{_zz_COMB_CSR__37,{_zz_COMB_CSR__38,_zz_COMB_CSR__39}}}}}}};
  assign _zz_COMB_CSR__35 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__36 = 12'hb0e;
  assign _zz_COMB_CSR__37 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h32d);
  assign _zz_COMB_CSR__38 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb8d);
  assign _zz_COMB_CSR__39 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb0d),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h32c),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb8c),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb0c),{(_zz_COMB_CSR__40 == _zz_COMB_CSR__41),{_zz_COMB_CSR__42,{_zz_COMB_CSR__43,_zz_COMB_CSR__44}}}}}}};
  assign _zz_COMB_CSR__40 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__41 = 12'h32b;
  assign _zz_COMB_CSR__42 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb8b);
  assign _zz_COMB_CSR__43 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb0b);
  assign _zz_COMB_CSR__44 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h32a),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb8a),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb0a),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h329),{(_zz_COMB_CSR__45 == _zz_COMB_CSR__46),{_zz_COMB_CSR__47,{_zz_COMB_CSR__48,_zz_COMB_CSR__49}}}}}}};
  assign _zz_COMB_CSR__45 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__46 = 12'hb89;
  assign _zz_COMB_CSR__47 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb09);
  assign _zz_COMB_CSR__48 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h328);
  assign _zz_COMB_CSR__49 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb88),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb08),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h327),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb87),{(_zz_COMB_CSR__50 == _zz_COMB_CSR__51),{_zz_COMB_CSR__52,{_zz_COMB_CSR__53,_zz_COMB_CSR__54}}}}}}};
  assign _zz_COMB_CSR__50 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__51 = 12'hb07;
  assign _zz_COMB_CSR__52 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h326);
  assign _zz_COMB_CSR__53 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb86);
  assign _zz_COMB_CSR__54 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb06),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h325),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb85),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb05),{(_zz_COMB_CSR__55 == _zz_COMB_CSR__56),{_zz_COMB_CSR__57,{_zz_COMB_CSR__58,_zz_COMB_CSR__59}}}}}}};
  assign _zz_COMB_CSR__55 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR__56 = 12'h324;
  assign _zz_COMB_CSR__57 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb84);
  assign _zz_COMB_CSR__58 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb04);
  assign _zz_COMB_CSR__59 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h323),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb83),(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb03)}};
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_1 = 12'hc82;
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_2 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc80);
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_3 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc06);
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_4 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc05),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc04),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc03),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc02),{(_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_5 == _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_6),{_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_7,{_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_8,_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_9}}}}}}};
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_5 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_6 = 12'hc00;
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_7 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb86);
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_8 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb85);
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_9 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb84),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb83),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb82),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb80),{(_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_10 == _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_11),{_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_12,{_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_13,_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_14}}}}}}};
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_10 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_11 = 12'hb06;
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_12 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb05);
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_13 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb04);
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_14 = {(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb03),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb02),(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb00)}};
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented = COMB_CSR_324;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_1 = {COMB_CSR_260,{COMB_CSR_256,{COMB_CSR_322,{COMB_CSR_320,{COMB_CSR_321,{COMB_CSR_323,{COMB_CSR_261,{COMB_CSR_771,{COMB_CSR_770,{COMB_CSR_772,{_zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_2,_zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_3}}}}}}}}}}};
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_2 = COMB_CSR_836;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_3 = {COMB_CSR_768,{COMB_CSR_834,{COMB_CSR_769,{COMB_CSR_3860,{COMB_CSR_3859,{COMB_CSR_3858,{COMB_CSR_3857,{COMB_CSR_832,{COMB_CSR_833,{COMB_CSR_835,COMB_CSR_773}}}}}}}}}};
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 = (REG_CSR_3857 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 = (REG_CSR_3858 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23 = (REG_CSR_3859 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 = (REG_CSR_3860 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29 = (REG_CSR_769 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31 = (REG_CSR_834 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33 = (REG_CSR_768 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35 = (REG_CSR_836 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37 = (REG_CSR_772 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39 = (REG_CSR_770 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41 = (REG_CSR_771 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43 = (REG_CSR_322 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45 = (REG_CSR_256 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47 = (REG_CSR_260 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49 = (REG_CSR_324 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51 = (REG_CSR_803 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50 = 32'h00000000;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52 = 32'h00000000;
  assign _zz_FrontendPlugin_decoded_LEGAL_0 = 32'h0000107f;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_1 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000207f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_2 = 32'h00002073;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_3 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000407f) == 32'h00004063);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_4 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000207f) == 32'h00002013);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_5 = {((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000107f) == 32'h00000013),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000603f) == 32'h00000023),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_LEGAL_0_6) == 32'h00000003),{(_zz_FrontendPlugin_decoded_LEGAL_0_7 == _zz_FrontendPlugin_decoded_LEGAL_0_8),{_zz_FrontendPlugin_decoded_LEGAL_0_9,{_zz_FrontendPlugin_decoded_LEGAL_0_10,_zz_FrontendPlugin_decoded_LEGAL_0_11}}}}}};
  assign _zz_FrontendPlugin_decoded_LEGAL_0_6 = 32'h0000207f;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_7 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000505f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_8 = 32'h00000003;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_9 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000707b) == 32'h00000063);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_10 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000607f) == 32'h0000000f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_11 = {((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h1800707f) == 32'h0000202f),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hfc00007f) == 32'h00000033),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_LEGAL_0_12) == 32'h0800202f),{(_zz_FrontendPlugin_decoded_LEGAL_0_13 == _zz_FrontendPlugin_decoded_LEGAL_0_14),{_zz_FrontendPlugin_decoded_LEGAL_0_15,{_zz_FrontendPlugin_decoded_LEGAL_0_16,_zz_FrontendPlugin_decoded_LEGAL_0_17}}}}}};
  assign _zz_FrontendPlugin_decoded_LEGAL_0_12 = 32'he800707f;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_13 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hfc00305f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_14 = 32'h00001013;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_15 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h01f0707f) == 32'h0000500f);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_16 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hbc00707f) == 32'h00005013);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_17 = {((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hbe00707f) == 32'h00005033),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hbe00707f) == 32'h00000033),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_LEGAL_0_18) == 32'h1000202f),{(_zz_FrontendPlugin_decoded_LEGAL_0_19 == _zz_FrontendPlugin_decoded_LEGAL_0_20),{_zz_FrontendPlugin_decoded_LEGAL_0_21,{_zz_FrontendPlugin_decoded_LEGAL_0_22,_zz_FrontendPlugin_decoded_LEGAL_0_23}}}}}};
  assign _zz_FrontendPlugin_decoded_LEGAL_0_18 = 32'hf9f0707f;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_19 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hfe007fff);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_20 = 32'h12000073;
  assign _zz_FrontendPlugin_decoded_LEGAL_0_21 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hdfffffff) == 32'h10200073);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_22 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hffefffff) == 32'h00000073);
  assign _zz_FrontendPlugin_decoded_LEGAL_0_23 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'hffffffff) == 32'h10500073);
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_2 = 32'h00002008;
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_3 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000050);
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_4 = 32'h00000010;
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0_5 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000028) == 32'h00000000);
  assign _zz_FrontendPlugin_decoded_LEGAL_1 = 32'h0000107f;
  assign _zz_FrontendPlugin_decoded_LEGAL_1_1 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000207f);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_2 = 32'h00002073;
  assign _zz_FrontendPlugin_decoded_LEGAL_1_3 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000407f) == 32'h00004063);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_4 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000207f) == 32'h00002013);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_5 = {((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000107f) == 32'h00000013),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000603f) == 32'h00000023),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & _zz_FrontendPlugin_decoded_LEGAL_1_6) == 32'h00000003),{(_zz_FrontendPlugin_decoded_LEGAL_1_7 == _zz_FrontendPlugin_decoded_LEGAL_1_8),{_zz_FrontendPlugin_decoded_LEGAL_1_9,{_zz_FrontendPlugin_decoded_LEGAL_1_10,_zz_FrontendPlugin_decoded_LEGAL_1_11}}}}}};
  assign _zz_FrontendPlugin_decoded_LEGAL_1_6 = 32'h0000207f;
  assign _zz_FrontendPlugin_decoded_LEGAL_1_7 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000505f);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_8 = 32'h00000003;
  assign _zz_FrontendPlugin_decoded_LEGAL_1_9 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000707b) == 32'h00000063);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_10 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000607f) == 32'h0000000f);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_11 = {((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h1800707f) == 32'h0000202f),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'hfc00007f) == 32'h00000033),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & _zz_FrontendPlugin_decoded_LEGAL_1_12) == 32'h0800202f),{(_zz_FrontendPlugin_decoded_LEGAL_1_13 == _zz_FrontendPlugin_decoded_LEGAL_1_14),{_zz_FrontendPlugin_decoded_LEGAL_1_15,{_zz_FrontendPlugin_decoded_LEGAL_1_16,_zz_FrontendPlugin_decoded_LEGAL_1_17}}}}}};
  assign _zz_FrontendPlugin_decoded_LEGAL_1_12 = 32'he800707f;
  assign _zz_FrontendPlugin_decoded_LEGAL_1_13 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'hfc00305f);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_14 = 32'h00001013;
  assign _zz_FrontendPlugin_decoded_LEGAL_1_15 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h01f0707f) == 32'h0000500f);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_16 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'hbc00707f) == 32'h00005013);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_17 = {((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'hbe00707f) == 32'h00005033),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'hbe00707f) == 32'h00000033),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & _zz_FrontendPlugin_decoded_LEGAL_1_18) == 32'h1000202f),{(_zz_FrontendPlugin_decoded_LEGAL_1_19 == _zz_FrontendPlugin_decoded_LEGAL_1_20),{_zz_FrontendPlugin_decoded_LEGAL_1_21,{_zz_FrontendPlugin_decoded_LEGAL_1_22,_zz_FrontendPlugin_decoded_LEGAL_1_23}}}}}};
  assign _zz_FrontendPlugin_decoded_LEGAL_1_18 = 32'hf9f0707f;
  assign _zz_FrontendPlugin_decoded_LEGAL_1_19 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'hfe007fff);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_20 = 32'h12000073;
  assign _zz_FrontendPlugin_decoded_LEGAL_1_21 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'hdfffffff) == 32'h10200073);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_22 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'hffefffff) == 32'h00000073);
  assign _zz_FrontendPlugin_decoded_LEGAL_1_23 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'hffffffff) == 32'h10500073);
  assign _zz_FrontendPlugin_decoded_WRITE_RD_1_1 = 32'h00002008;
  assign _zz_FrontendPlugin_decoded_WRITE_RD_1_2 = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000050);
  assign _zz_FrontendPlugin_decoded_WRITE_RD_1_3 = 32'h00000010;
  assign _zz_FrontendPlugin_decoded_WRITE_RD_1_4 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000028) == 32'h00000000);
  assign _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0 = DispatchPlugin_logic_queue_io_contexts_24_staticWake[0];
  assign _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_1 = DispatchPlugin_logic_queue_io_contexts_23_staticWake[0];
  assign _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_2 = {DispatchPlugin_logic_queue_io_contexts_22_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_21_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_20_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_19_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_18_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_17_staticWake[0],{_zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_3,{_zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_4,_zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_5}}}}}}}};
  assign _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_3 = DispatchPlugin_logic_queue_io_contexts_16_staticWake[0];
  assign _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_4 = DispatchPlugin_logic_queue_io_contexts_15_staticWake[0];
  assign _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_5 = {DispatchPlugin_logic_queue_io_contexts_14_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_13_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_12_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_11_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_10_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_9_staticWake[0],{_zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_6,{_zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_7,_zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_8}}}}}}}};
  assign _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_6 = DispatchPlugin_logic_queue_io_contexts_8_staticWake[0];
  assign _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_7 = DispatchPlugin_logic_queue_io_contexts_7_staticWake[0];
  assign _zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_8 = {DispatchPlugin_logic_queue_io_contexts_6_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_5_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_4_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_3_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_2_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_1_staticWake[0],DispatchPlugin_logic_queue_io_contexts_0_staticWake[0]}}}}}};
  assign _zz_DispatchPlugin_logic_pop_0_portEventFull = 1'b0;
  assign _zz_DispatchPlugin_logic_pop_0_portEventFull_1 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[11];
  assign _zz_DispatchPlugin_logic_pop_0_portEventFull_2 = {1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[10],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[9],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[8],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[7],{1'b0,{_zz_DispatchPlugin_logic_pop_0_portEventFull_3,{_zz_DispatchPlugin_logic_pop_0_portEventFull_4,_zz_DispatchPlugin_logic_pop_0_portEventFull_5}}}}}}}}}}};
  assign _zz_DispatchPlugin_logic_pop_0_portEventFull_3 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[6];
  assign _zz_DispatchPlugin_logic_pop_0_portEventFull_4 = 1'b0;
  assign _zz_DispatchPlugin_logic_pop_0_portEventFull_5 = {DispatchPlugin_logic_queue_io_schedules_0_payload_event[5],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[4],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[3],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[2],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[1],{_zz_DispatchPlugin_logic_pop_0_portEventFull_6,_zz_DispatchPlugin_logic_pop_0_portEventFull_7}}}}}}}}}};
  assign _zz_DispatchPlugin_logic_pop_0_portEventFull_6 = 1'b0;
  assign _zz_DispatchPlugin_logic_pop_0_portEventFull_7 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[0];
  assign _zz_DispatchPlugin_logic_pop_1_portEventFull = DispatchPlugin_logic_queue_io_schedules_1_payload_event[11];
  assign _zz_DispatchPlugin_logic_pop_1_portEventFull_1 = 1'b0;
  assign _zz_DispatchPlugin_logic_pop_1_portEventFull_2 = {DispatchPlugin_logic_queue_io_schedules_1_payload_event[10],{1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[9],{1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[8],{1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[7],{_zz_DispatchPlugin_logic_pop_1_portEventFull_3,{_zz_DispatchPlugin_logic_pop_1_portEventFull_4,_zz_DispatchPlugin_logic_pop_1_portEventFull_5}}}}}}}}};
  assign _zz_DispatchPlugin_logic_pop_1_portEventFull_3 = 1'b0;
  assign _zz_DispatchPlugin_logic_pop_1_portEventFull_4 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[6];
  assign _zz_DispatchPlugin_logic_pop_1_portEventFull_5 = {1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[5],{1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[4],{1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[3],{1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[2],{1'b0,{_zz_DispatchPlugin_logic_pop_1_portEventFull_6,{_zz_DispatchPlugin_logic_pop_1_portEventFull_7,_zz_DispatchPlugin_logic_pop_1_portEventFull_8}}}}}}}}}}};
  assign _zz_DispatchPlugin_logic_pop_1_portEventFull_6 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[1];
  assign _zz_DispatchPlugin_logic_pop_1_portEventFull_7 = 1'b0;
  assign _zz_DispatchPlugin_logic_pop_1_portEventFull_8 = {DispatchPlugin_logic_queue_io_schedules_1_payload_event[0],1'b0};
  assign _zz_DispatchPlugin_logic_pop_2_portEventFull = DispatchPlugin_logic_queue_io_schedules_2_payload_event[24];
  assign _zz_DispatchPlugin_logic_pop_2_portEventFull_1 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[23];
  assign _zz_DispatchPlugin_logic_pop_2_portEventFull_2 = {DispatchPlugin_logic_queue_io_schedules_2_payload_event[22],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[21],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[20],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[19],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[18],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[17],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[16],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[15],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[14],{_zz_DispatchPlugin_logic_pop_2_portEventFull_3,{_zz_DispatchPlugin_logic_pop_2_portEventFull_4,_zz_DispatchPlugin_logic_pop_2_portEventFull_5}}}}}}}}}}};
  assign _zz_DispatchPlugin_logic_pop_2_portEventFull_3 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[13];
  assign _zz_DispatchPlugin_logic_pop_2_portEventFull_4 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[12];
  assign _zz_DispatchPlugin_logic_pop_2_portEventFull_5 = {DispatchPlugin_logic_queue_io_schedules_2_payload_event[11],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[10],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[9],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[8],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[7],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[6],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[5],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[4],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[3],{_zz_DispatchPlugin_logic_pop_2_portEventFull_6,{_zz_DispatchPlugin_logic_pop_2_portEventFull_7,_zz_DispatchPlugin_logic_pop_2_portEventFull_8}}}}}}}}}}};
  assign _zz_DispatchPlugin_logic_pop_2_portEventFull_6 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[2];
  assign _zz_DispatchPlugin_logic_pop_2_portEventFull_7 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[1];
  assign _zz_DispatchPlugin_logic_pop_2_portEventFull_8 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[0];
  always @(posedge clk) begin
    if(_zz_when_MultiportRam_l328_4) begin
      FetchCachePlugin_logic_banks_0_mem[FetchCachePlugin_logic_banks_0_write_payload_address] <= FetchCachePlugin_logic_banks_0_write_payload_data;
    end
  end

  always @(posedge clk) begin
    if(FetchCachePlugin_logic_banks_0_read_cmd_valid) begin
      _zz_FetchCachePlugin_logic_banks_0_mem_port1 <= FetchCachePlugin_logic_banks_0_mem[FetchCachePlugin_logic_banks_0_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_when_MultiportRam_l328_3) begin
      FetchCachePlugin_logic_banks_1_mem[FetchCachePlugin_logic_banks_1_write_payload_address] <= FetchCachePlugin_logic_banks_1_write_payload_data;
    end
  end

  always @(posedge clk) begin
    if(FetchCachePlugin_logic_banks_1_read_cmd_valid) begin
      _zz_FetchCachePlugin_logic_banks_1_mem_port1 <= FetchCachePlugin_logic_banks_1_mem[FetchCachePlugin_logic_banks_1_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_when_MultiportRam_l328_2) begin
      FetchCachePlugin_logic_banks_2_mem[FetchCachePlugin_logic_banks_2_write_payload_address] <= FetchCachePlugin_logic_banks_2_write_payload_data;
    end
  end

  always @(posedge clk) begin
    if(FetchCachePlugin_logic_banks_2_read_cmd_valid) begin
      _zz_FetchCachePlugin_logic_banks_2_mem_port1 <= FetchCachePlugin_logic_banks_2_mem[FetchCachePlugin_logic_banks_2_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_when_MultiportRam_l328_1) begin
      FetchCachePlugin_logic_banks_3_mem[FetchCachePlugin_logic_banks_3_write_payload_address] <= FetchCachePlugin_logic_banks_3_write_payload_data;
    end
  end

  always @(posedge clk) begin
    if(FetchCachePlugin_logic_banks_3_read_cmd_valid) begin
      _zz_FetchCachePlugin_logic_banks_3_mem_port1 <= FetchCachePlugin_logic_banks_3_mem[FetchCachePlugin_logic_banks_3_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_logic_ways_0_mem_port_1) begin
      FetchCachePlugin_logic_ways_0_mem[FetchCachePlugin_logic_waysWrite_address] <= _zz_FetchCachePlugin_logic_ways_0_mem_port;
    end
  end

  assign _zz_FetchCachePlugin_logic_ways_0_mem_port1 = FetchCachePlugin_logic_ways_0_mem[FetchCachePlugin_logic_ways_0_read_cmd_payload];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_logic_ways_1_mem_port_1) begin
      FetchCachePlugin_logic_ways_1_mem[FetchCachePlugin_logic_waysWrite_address] <= _zz_FetchCachePlugin_logic_ways_1_mem_port;
    end
  end

  assign _zz_FetchCachePlugin_logic_ways_1_mem_port1 = FetchCachePlugin_logic_ways_1_mem[FetchCachePlugin_logic_ways_1_read_cmd_payload];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_logic_ways_2_mem_port_1) begin
      FetchCachePlugin_logic_ways_2_mem[FetchCachePlugin_logic_waysWrite_address] <= _zz_FetchCachePlugin_logic_ways_2_mem_port;
    end
  end

  assign _zz_FetchCachePlugin_logic_ways_2_mem_port1 = FetchCachePlugin_logic_ways_2_mem[FetchCachePlugin_logic_ways_2_read_cmd_payload];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_logic_ways_3_mem_port_1) begin
      FetchCachePlugin_logic_ways_3_mem[FetchCachePlugin_logic_waysWrite_address] <= _zz_FetchCachePlugin_logic_ways_3_mem_port;
    end
  end

  assign _zz_FetchCachePlugin_logic_ways_3_mem_port1 = FetchCachePlugin_logic_ways_3_mem[FetchCachePlugin_logic_ways_3_read_cmd_payload];
  always @(posedge clk) begin
    if(_zz_18) begin
      FetchCachePlugin_logic_plru_ram[FetchCachePlugin_logic_plru_write_payload_address] <= _zz_FetchCachePlugin_logic_plru_ram_port;
    end
  end

  assign _zz_FetchCachePlugin_logic_plru_ram_port1 = FetchCachePlugin_logic_plru_ram[_zz_FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0];
  initial begin
    DecoderPredictionPlugin_logic_ras_mem_stack[0] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[1] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[2] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[3] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[4] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[5] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[6] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[7] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[8] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[9] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[10] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[11] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[12] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[13] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[14] = 32'b00000000000000000000000000000000;
    DecoderPredictionPlugin_logic_ras_mem_stack[15] = 32'b00000000000000000000000000000000;
  end
  assign _zz_DecoderPredictionPlugin_logic_ras_mem_stack_port0 = DecoderPredictionPlugin_logic_ras_mem_stack[DecoderPredictionPlugin_logic_ras_ptr_pop];
  always @(posedge clk) begin
    if(_zz_17) begin
      DecoderPredictionPlugin_logic_ras_mem_stack[DecoderPredictionPlugin_logic_ras_write_payload_address] <= _zz_DecoderPredictionPlugin_logic_ras_mem_stack_port;
    end
  end

  initial begin
    BtbPlugin_logic_mem[0] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[1] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[2] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[3] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[4] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[5] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[6] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[7] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[8] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[9] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[10] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[11] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[12] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[13] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[14] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[15] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[16] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[17] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[18] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[19] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[20] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[21] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[22] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[23] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[24] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[25] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[26] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[27] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[28] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[29] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[30] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[31] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[32] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[33] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[34] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[35] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[36] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[37] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[38] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[39] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[40] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[41] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[42] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[43] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[44] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[45] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[46] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[47] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[48] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[49] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[50] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[51] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[52] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[53] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[54] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[55] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[56] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[57] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[58] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[59] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[60] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[61] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[62] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[63] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[64] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[65] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[66] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[67] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[68] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[69] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[70] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[71] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[72] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[73] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[74] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[75] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[76] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[77] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[78] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[79] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[80] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[81] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[82] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[83] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[84] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[85] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[86] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[87] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[88] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[89] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[90] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[91] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[92] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[93] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[94] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[95] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[96] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[97] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[98] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[99] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[100] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[101] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[102] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[103] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[104] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[105] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[106] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[107] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[108] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[109] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[110] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[111] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[112] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[113] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[114] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[115] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[116] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[117] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[118] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[119] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[120] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[121] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[122] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[123] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[124] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[125] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[126] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[127] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[128] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[129] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[130] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[131] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[132] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[133] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[134] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[135] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[136] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[137] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[138] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[139] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[140] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[141] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[142] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[143] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[144] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[145] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[146] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[147] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[148] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[149] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[150] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[151] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[152] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[153] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[154] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[155] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[156] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[157] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[158] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[159] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[160] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[161] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[162] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[163] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[164] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[165] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[166] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[167] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[168] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[169] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[170] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[171] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[172] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[173] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[174] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[175] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[176] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[177] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[178] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[179] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[180] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[181] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[182] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[183] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[184] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[185] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[186] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[187] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[188] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[189] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[190] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[191] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[192] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[193] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[194] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[195] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[196] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[197] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[198] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[199] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[200] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[201] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[202] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[203] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[204] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[205] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[206] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[207] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[208] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[209] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[210] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[211] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[212] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[213] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[214] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[215] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[216] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[217] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[218] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[219] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[220] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[221] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[222] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[223] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[224] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[225] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[226] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[227] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[228] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[229] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[230] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[231] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[232] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[233] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[234] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[235] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[236] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[237] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[238] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[239] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[240] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[241] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[242] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[243] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[244] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[245] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[246] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[247] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[248] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[249] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[250] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[251] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[252] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[253] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[254] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[255] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[256] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[257] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[258] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[259] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[260] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[261] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[262] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[263] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[264] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[265] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[266] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[267] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[268] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[269] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[270] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[271] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[272] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[273] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[274] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[275] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[276] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[277] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[278] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[279] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[280] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[281] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[282] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[283] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[284] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[285] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[286] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[287] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[288] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[289] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[290] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[291] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[292] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[293] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[294] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[295] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[296] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[297] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[298] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[299] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[300] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[301] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[302] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[303] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[304] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[305] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[306] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[307] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[308] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[309] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[310] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[311] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[312] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[313] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[314] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[315] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[316] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[317] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[318] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[319] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[320] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[321] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[322] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[323] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[324] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[325] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[326] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[327] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[328] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[329] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[330] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[331] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[332] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[333] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[334] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[335] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[336] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[337] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[338] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[339] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[340] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[341] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[342] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[343] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[344] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[345] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[346] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[347] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[348] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[349] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[350] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[351] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[352] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[353] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[354] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[355] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[356] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[357] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[358] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[359] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[360] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[361] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[362] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[363] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[364] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[365] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[366] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[367] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[368] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[369] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[370] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[371] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[372] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[373] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[374] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[375] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[376] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[377] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[378] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[379] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[380] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[381] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[382] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[383] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[384] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[385] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[386] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[387] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[388] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[389] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[390] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[391] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[392] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[393] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[394] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[395] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[396] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[397] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[398] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[399] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[400] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[401] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[402] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[403] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[404] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[405] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[406] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[407] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[408] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[409] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[410] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[411] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[412] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[413] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[414] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[415] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[416] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[417] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[418] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[419] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[420] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[421] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[422] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[423] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[424] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[425] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[426] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[427] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[428] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[429] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[430] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[431] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[432] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[433] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[434] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[435] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[436] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[437] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[438] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[439] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[440] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[441] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[442] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[443] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[444] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[445] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[446] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[447] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[448] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[449] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[450] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[451] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[452] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[453] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[454] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[455] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[456] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[457] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[458] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[459] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[460] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[461] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[462] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[463] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[464] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[465] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[466] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[467] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[468] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[469] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[470] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[471] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[472] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[473] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[474] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[475] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[476] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[477] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[478] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[479] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[480] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[481] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[482] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[483] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[484] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[485] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[486] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[487] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[488] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[489] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[490] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[491] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[492] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[493] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[494] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[495] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[496] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[497] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[498] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[499] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[500] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[501] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[502] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[503] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[504] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[505] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[506] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[507] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[508] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[509] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[510] = 50'b00000000000000000000000000000000000000000000000000;
    BtbPlugin_logic_mem[511] = 50'b00000000000000000000000000000000000000000000000000;
  end
  always @(posedge clk) begin
    if(FetchPlugin_stages_0_ready) begin
      _zz_BtbPlugin_logic_mem_port1 <= BtbPlugin_logic_mem[BtbPlugin_logic_readCmd_entryAddress];
    end
    if(_zz_16) begin
      BtbPlugin_logic_mem[BtbPlugin_logic_onLearn_port_payload_address] <= _zz_BtbPlugin_logic_mem_port;
    end
  end

  initial begin
    GSharePlugin_logic_mem_counter[0] = 4'b0000;
    GSharePlugin_logic_mem_counter[1] = 4'b0000;
    GSharePlugin_logic_mem_counter[2] = 4'b0000;
    GSharePlugin_logic_mem_counter[3] = 4'b0000;
    GSharePlugin_logic_mem_counter[4] = 4'b0000;
    GSharePlugin_logic_mem_counter[5] = 4'b0000;
    GSharePlugin_logic_mem_counter[6] = 4'b0000;
    GSharePlugin_logic_mem_counter[7] = 4'b0000;
    GSharePlugin_logic_mem_counter[8] = 4'b0000;
    GSharePlugin_logic_mem_counter[9] = 4'b0000;
    GSharePlugin_logic_mem_counter[10] = 4'b0000;
    GSharePlugin_logic_mem_counter[11] = 4'b0000;
    GSharePlugin_logic_mem_counter[12] = 4'b0000;
    GSharePlugin_logic_mem_counter[13] = 4'b0000;
    GSharePlugin_logic_mem_counter[14] = 4'b0000;
    GSharePlugin_logic_mem_counter[15] = 4'b0000;
    GSharePlugin_logic_mem_counter[16] = 4'b0000;
    GSharePlugin_logic_mem_counter[17] = 4'b0000;
    GSharePlugin_logic_mem_counter[18] = 4'b0000;
    GSharePlugin_logic_mem_counter[19] = 4'b0000;
    GSharePlugin_logic_mem_counter[20] = 4'b0000;
    GSharePlugin_logic_mem_counter[21] = 4'b0000;
    GSharePlugin_logic_mem_counter[22] = 4'b0000;
    GSharePlugin_logic_mem_counter[23] = 4'b0000;
    GSharePlugin_logic_mem_counter[24] = 4'b0000;
    GSharePlugin_logic_mem_counter[25] = 4'b0000;
    GSharePlugin_logic_mem_counter[26] = 4'b0000;
    GSharePlugin_logic_mem_counter[27] = 4'b0000;
    GSharePlugin_logic_mem_counter[28] = 4'b0000;
    GSharePlugin_logic_mem_counter[29] = 4'b0000;
    GSharePlugin_logic_mem_counter[30] = 4'b0000;
    GSharePlugin_logic_mem_counter[31] = 4'b0000;
    GSharePlugin_logic_mem_counter[32] = 4'b0000;
    GSharePlugin_logic_mem_counter[33] = 4'b0000;
    GSharePlugin_logic_mem_counter[34] = 4'b0000;
    GSharePlugin_logic_mem_counter[35] = 4'b0000;
    GSharePlugin_logic_mem_counter[36] = 4'b0000;
    GSharePlugin_logic_mem_counter[37] = 4'b0000;
    GSharePlugin_logic_mem_counter[38] = 4'b0000;
    GSharePlugin_logic_mem_counter[39] = 4'b0000;
    GSharePlugin_logic_mem_counter[40] = 4'b0000;
    GSharePlugin_logic_mem_counter[41] = 4'b0000;
    GSharePlugin_logic_mem_counter[42] = 4'b0000;
    GSharePlugin_logic_mem_counter[43] = 4'b0000;
    GSharePlugin_logic_mem_counter[44] = 4'b0000;
    GSharePlugin_logic_mem_counter[45] = 4'b0000;
    GSharePlugin_logic_mem_counter[46] = 4'b0000;
    GSharePlugin_logic_mem_counter[47] = 4'b0000;
    GSharePlugin_logic_mem_counter[48] = 4'b0000;
    GSharePlugin_logic_mem_counter[49] = 4'b0000;
    GSharePlugin_logic_mem_counter[50] = 4'b0000;
    GSharePlugin_logic_mem_counter[51] = 4'b0000;
    GSharePlugin_logic_mem_counter[52] = 4'b0000;
    GSharePlugin_logic_mem_counter[53] = 4'b0000;
    GSharePlugin_logic_mem_counter[54] = 4'b0000;
    GSharePlugin_logic_mem_counter[55] = 4'b0000;
    GSharePlugin_logic_mem_counter[56] = 4'b0000;
    GSharePlugin_logic_mem_counter[57] = 4'b0000;
    GSharePlugin_logic_mem_counter[58] = 4'b0000;
    GSharePlugin_logic_mem_counter[59] = 4'b0000;
    GSharePlugin_logic_mem_counter[60] = 4'b0000;
    GSharePlugin_logic_mem_counter[61] = 4'b0000;
    GSharePlugin_logic_mem_counter[62] = 4'b0000;
    GSharePlugin_logic_mem_counter[63] = 4'b0000;
    GSharePlugin_logic_mem_counter[64] = 4'b0000;
    GSharePlugin_logic_mem_counter[65] = 4'b0000;
    GSharePlugin_logic_mem_counter[66] = 4'b0000;
    GSharePlugin_logic_mem_counter[67] = 4'b0000;
    GSharePlugin_logic_mem_counter[68] = 4'b0000;
    GSharePlugin_logic_mem_counter[69] = 4'b0000;
    GSharePlugin_logic_mem_counter[70] = 4'b0000;
    GSharePlugin_logic_mem_counter[71] = 4'b0000;
    GSharePlugin_logic_mem_counter[72] = 4'b0000;
    GSharePlugin_logic_mem_counter[73] = 4'b0000;
    GSharePlugin_logic_mem_counter[74] = 4'b0000;
    GSharePlugin_logic_mem_counter[75] = 4'b0000;
    GSharePlugin_logic_mem_counter[76] = 4'b0000;
    GSharePlugin_logic_mem_counter[77] = 4'b0000;
    GSharePlugin_logic_mem_counter[78] = 4'b0000;
    GSharePlugin_logic_mem_counter[79] = 4'b0000;
    GSharePlugin_logic_mem_counter[80] = 4'b0000;
    GSharePlugin_logic_mem_counter[81] = 4'b0000;
    GSharePlugin_logic_mem_counter[82] = 4'b0000;
    GSharePlugin_logic_mem_counter[83] = 4'b0000;
    GSharePlugin_logic_mem_counter[84] = 4'b0000;
    GSharePlugin_logic_mem_counter[85] = 4'b0000;
    GSharePlugin_logic_mem_counter[86] = 4'b0000;
    GSharePlugin_logic_mem_counter[87] = 4'b0000;
    GSharePlugin_logic_mem_counter[88] = 4'b0000;
    GSharePlugin_logic_mem_counter[89] = 4'b0000;
    GSharePlugin_logic_mem_counter[90] = 4'b0000;
    GSharePlugin_logic_mem_counter[91] = 4'b0000;
    GSharePlugin_logic_mem_counter[92] = 4'b0000;
    GSharePlugin_logic_mem_counter[93] = 4'b0000;
    GSharePlugin_logic_mem_counter[94] = 4'b0000;
    GSharePlugin_logic_mem_counter[95] = 4'b0000;
    GSharePlugin_logic_mem_counter[96] = 4'b0000;
    GSharePlugin_logic_mem_counter[97] = 4'b0000;
    GSharePlugin_logic_mem_counter[98] = 4'b0000;
    GSharePlugin_logic_mem_counter[99] = 4'b0000;
    GSharePlugin_logic_mem_counter[100] = 4'b0000;
    GSharePlugin_logic_mem_counter[101] = 4'b0000;
    GSharePlugin_logic_mem_counter[102] = 4'b0000;
    GSharePlugin_logic_mem_counter[103] = 4'b0000;
    GSharePlugin_logic_mem_counter[104] = 4'b0000;
    GSharePlugin_logic_mem_counter[105] = 4'b0000;
    GSharePlugin_logic_mem_counter[106] = 4'b0000;
    GSharePlugin_logic_mem_counter[107] = 4'b0000;
    GSharePlugin_logic_mem_counter[108] = 4'b0000;
    GSharePlugin_logic_mem_counter[109] = 4'b0000;
    GSharePlugin_logic_mem_counter[110] = 4'b0000;
    GSharePlugin_logic_mem_counter[111] = 4'b0000;
    GSharePlugin_logic_mem_counter[112] = 4'b0000;
    GSharePlugin_logic_mem_counter[113] = 4'b0000;
    GSharePlugin_logic_mem_counter[114] = 4'b0000;
    GSharePlugin_logic_mem_counter[115] = 4'b0000;
    GSharePlugin_logic_mem_counter[116] = 4'b0000;
    GSharePlugin_logic_mem_counter[117] = 4'b0000;
    GSharePlugin_logic_mem_counter[118] = 4'b0000;
    GSharePlugin_logic_mem_counter[119] = 4'b0000;
    GSharePlugin_logic_mem_counter[120] = 4'b0000;
    GSharePlugin_logic_mem_counter[121] = 4'b0000;
    GSharePlugin_logic_mem_counter[122] = 4'b0000;
    GSharePlugin_logic_mem_counter[123] = 4'b0000;
    GSharePlugin_logic_mem_counter[124] = 4'b0000;
    GSharePlugin_logic_mem_counter[125] = 4'b0000;
    GSharePlugin_logic_mem_counter[126] = 4'b0000;
    GSharePlugin_logic_mem_counter[127] = 4'b0000;
    GSharePlugin_logic_mem_counter[128] = 4'b0000;
    GSharePlugin_logic_mem_counter[129] = 4'b0000;
    GSharePlugin_logic_mem_counter[130] = 4'b0000;
    GSharePlugin_logic_mem_counter[131] = 4'b0000;
    GSharePlugin_logic_mem_counter[132] = 4'b0000;
    GSharePlugin_logic_mem_counter[133] = 4'b0000;
    GSharePlugin_logic_mem_counter[134] = 4'b0000;
    GSharePlugin_logic_mem_counter[135] = 4'b0000;
    GSharePlugin_logic_mem_counter[136] = 4'b0000;
    GSharePlugin_logic_mem_counter[137] = 4'b0000;
    GSharePlugin_logic_mem_counter[138] = 4'b0000;
    GSharePlugin_logic_mem_counter[139] = 4'b0000;
    GSharePlugin_logic_mem_counter[140] = 4'b0000;
    GSharePlugin_logic_mem_counter[141] = 4'b0000;
    GSharePlugin_logic_mem_counter[142] = 4'b0000;
    GSharePlugin_logic_mem_counter[143] = 4'b0000;
    GSharePlugin_logic_mem_counter[144] = 4'b0000;
    GSharePlugin_logic_mem_counter[145] = 4'b0000;
    GSharePlugin_logic_mem_counter[146] = 4'b0000;
    GSharePlugin_logic_mem_counter[147] = 4'b0000;
    GSharePlugin_logic_mem_counter[148] = 4'b0000;
    GSharePlugin_logic_mem_counter[149] = 4'b0000;
    GSharePlugin_logic_mem_counter[150] = 4'b0000;
    GSharePlugin_logic_mem_counter[151] = 4'b0000;
    GSharePlugin_logic_mem_counter[152] = 4'b0000;
    GSharePlugin_logic_mem_counter[153] = 4'b0000;
    GSharePlugin_logic_mem_counter[154] = 4'b0000;
    GSharePlugin_logic_mem_counter[155] = 4'b0000;
    GSharePlugin_logic_mem_counter[156] = 4'b0000;
    GSharePlugin_logic_mem_counter[157] = 4'b0000;
    GSharePlugin_logic_mem_counter[158] = 4'b0000;
    GSharePlugin_logic_mem_counter[159] = 4'b0000;
    GSharePlugin_logic_mem_counter[160] = 4'b0000;
    GSharePlugin_logic_mem_counter[161] = 4'b0000;
    GSharePlugin_logic_mem_counter[162] = 4'b0000;
    GSharePlugin_logic_mem_counter[163] = 4'b0000;
    GSharePlugin_logic_mem_counter[164] = 4'b0000;
    GSharePlugin_logic_mem_counter[165] = 4'b0000;
    GSharePlugin_logic_mem_counter[166] = 4'b0000;
    GSharePlugin_logic_mem_counter[167] = 4'b0000;
    GSharePlugin_logic_mem_counter[168] = 4'b0000;
    GSharePlugin_logic_mem_counter[169] = 4'b0000;
    GSharePlugin_logic_mem_counter[170] = 4'b0000;
    GSharePlugin_logic_mem_counter[171] = 4'b0000;
    GSharePlugin_logic_mem_counter[172] = 4'b0000;
    GSharePlugin_logic_mem_counter[173] = 4'b0000;
    GSharePlugin_logic_mem_counter[174] = 4'b0000;
    GSharePlugin_logic_mem_counter[175] = 4'b0000;
    GSharePlugin_logic_mem_counter[176] = 4'b0000;
    GSharePlugin_logic_mem_counter[177] = 4'b0000;
    GSharePlugin_logic_mem_counter[178] = 4'b0000;
    GSharePlugin_logic_mem_counter[179] = 4'b0000;
    GSharePlugin_logic_mem_counter[180] = 4'b0000;
    GSharePlugin_logic_mem_counter[181] = 4'b0000;
    GSharePlugin_logic_mem_counter[182] = 4'b0000;
    GSharePlugin_logic_mem_counter[183] = 4'b0000;
    GSharePlugin_logic_mem_counter[184] = 4'b0000;
    GSharePlugin_logic_mem_counter[185] = 4'b0000;
    GSharePlugin_logic_mem_counter[186] = 4'b0000;
    GSharePlugin_logic_mem_counter[187] = 4'b0000;
    GSharePlugin_logic_mem_counter[188] = 4'b0000;
    GSharePlugin_logic_mem_counter[189] = 4'b0000;
    GSharePlugin_logic_mem_counter[190] = 4'b0000;
    GSharePlugin_logic_mem_counter[191] = 4'b0000;
    GSharePlugin_logic_mem_counter[192] = 4'b0000;
    GSharePlugin_logic_mem_counter[193] = 4'b0000;
    GSharePlugin_logic_mem_counter[194] = 4'b0000;
    GSharePlugin_logic_mem_counter[195] = 4'b0000;
    GSharePlugin_logic_mem_counter[196] = 4'b0000;
    GSharePlugin_logic_mem_counter[197] = 4'b0000;
    GSharePlugin_logic_mem_counter[198] = 4'b0000;
    GSharePlugin_logic_mem_counter[199] = 4'b0000;
    GSharePlugin_logic_mem_counter[200] = 4'b0000;
    GSharePlugin_logic_mem_counter[201] = 4'b0000;
    GSharePlugin_logic_mem_counter[202] = 4'b0000;
    GSharePlugin_logic_mem_counter[203] = 4'b0000;
    GSharePlugin_logic_mem_counter[204] = 4'b0000;
    GSharePlugin_logic_mem_counter[205] = 4'b0000;
    GSharePlugin_logic_mem_counter[206] = 4'b0000;
    GSharePlugin_logic_mem_counter[207] = 4'b0000;
    GSharePlugin_logic_mem_counter[208] = 4'b0000;
    GSharePlugin_logic_mem_counter[209] = 4'b0000;
    GSharePlugin_logic_mem_counter[210] = 4'b0000;
    GSharePlugin_logic_mem_counter[211] = 4'b0000;
    GSharePlugin_logic_mem_counter[212] = 4'b0000;
    GSharePlugin_logic_mem_counter[213] = 4'b0000;
    GSharePlugin_logic_mem_counter[214] = 4'b0000;
    GSharePlugin_logic_mem_counter[215] = 4'b0000;
    GSharePlugin_logic_mem_counter[216] = 4'b0000;
    GSharePlugin_logic_mem_counter[217] = 4'b0000;
    GSharePlugin_logic_mem_counter[218] = 4'b0000;
    GSharePlugin_logic_mem_counter[219] = 4'b0000;
    GSharePlugin_logic_mem_counter[220] = 4'b0000;
    GSharePlugin_logic_mem_counter[221] = 4'b0000;
    GSharePlugin_logic_mem_counter[222] = 4'b0000;
    GSharePlugin_logic_mem_counter[223] = 4'b0000;
    GSharePlugin_logic_mem_counter[224] = 4'b0000;
    GSharePlugin_logic_mem_counter[225] = 4'b0000;
    GSharePlugin_logic_mem_counter[226] = 4'b0000;
    GSharePlugin_logic_mem_counter[227] = 4'b0000;
    GSharePlugin_logic_mem_counter[228] = 4'b0000;
    GSharePlugin_logic_mem_counter[229] = 4'b0000;
    GSharePlugin_logic_mem_counter[230] = 4'b0000;
    GSharePlugin_logic_mem_counter[231] = 4'b0000;
    GSharePlugin_logic_mem_counter[232] = 4'b0000;
    GSharePlugin_logic_mem_counter[233] = 4'b0000;
    GSharePlugin_logic_mem_counter[234] = 4'b0000;
    GSharePlugin_logic_mem_counter[235] = 4'b0000;
    GSharePlugin_logic_mem_counter[236] = 4'b0000;
    GSharePlugin_logic_mem_counter[237] = 4'b0000;
    GSharePlugin_logic_mem_counter[238] = 4'b0000;
    GSharePlugin_logic_mem_counter[239] = 4'b0000;
    GSharePlugin_logic_mem_counter[240] = 4'b0000;
    GSharePlugin_logic_mem_counter[241] = 4'b0000;
    GSharePlugin_logic_mem_counter[242] = 4'b0000;
    GSharePlugin_logic_mem_counter[243] = 4'b0000;
    GSharePlugin_logic_mem_counter[244] = 4'b0000;
    GSharePlugin_logic_mem_counter[245] = 4'b0000;
    GSharePlugin_logic_mem_counter[246] = 4'b0000;
    GSharePlugin_logic_mem_counter[247] = 4'b0000;
    GSharePlugin_logic_mem_counter[248] = 4'b0000;
    GSharePlugin_logic_mem_counter[249] = 4'b0000;
    GSharePlugin_logic_mem_counter[250] = 4'b0000;
    GSharePlugin_logic_mem_counter[251] = 4'b0000;
    GSharePlugin_logic_mem_counter[252] = 4'b0000;
    GSharePlugin_logic_mem_counter[253] = 4'b0000;
    GSharePlugin_logic_mem_counter[254] = 4'b0000;
    GSharePlugin_logic_mem_counter[255] = 4'b0000;
    GSharePlugin_logic_mem_counter[256] = 4'b0000;
    GSharePlugin_logic_mem_counter[257] = 4'b0000;
    GSharePlugin_logic_mem_counter[258] = 4'b0000;
    GSharePlugin_logic_mem_counter[259] = 4'b0000;
    GSharePlugin_logic_mem_counter[260] = 4'b0000;
    GSharePlugin_logic_mem_counter[261] = 4'b0000;
    GSharePlugin_logic_mem_counter[262] = 4'b0000;
    GSharePlugin_logic_mem_counter[263] = 4'b0000;
    GSharePlugin_logic_mem_counter[264] = 4'b0000;
    GSharePlugin_logic_mem_counter[265] = 4'b0000;
    GSharePlugin_logic_mem_counter[266] = 4'b0000;
    GSharePlugin_logic_mem_counter[267] = 4'b0000;
    GSharePlugin_logic_mem_counter[268] = 4'b0000;
    GSharePlugin_logic_mem_counter[269] = 4'b0000;
    GSharePlugin_logic_mem_counter[270] = 4'b0000;
    GSharePlugin_logic_mem_counter[271] = 4'b0000;
    GSharePlugin_logic_mem_counter[272] = 4'b0000;
    GSharePlugin_logic_mem_counter[273] = 4'b0000;
    GSharePlugin_logic_mem_counter[274] = 4'b0000;
    GSharePlugin_logic_mem_counter[275] = 4'b0000;
    GSharePlugin_logic_mem_counter[276] = 4'b0000;
    GSharePlugin_logic_mem_counter[277] = 4'b0000;
    GSharePlugin_logic_mem_counter[278] = 4'b0000;
    GSharePlugin_logic_mem_counter[279] = 4'b0000;
    GSharePlugin_logic_mem_counter[280] = 4'b0000;
    GSharePlugin_logic_mem_counter[281] = 4'b0000;
    GSharePlugin_logic_mem_counter[282] = 4'b0000;
    GSharePlugin_logic_mem_counter[283] = 4'b0000;
    GSharePlugin_logic_mem_counter[284] = 4'b0000;
    GSharePlugin_logic_mem_counter[285] = 4'b0000;
    GSharePlugin_logic_mem_counter[286] = 4'b0000;
    GSharePlugin_logic_mem_counter[287] = 4'b0000;
    GSharePlugin_logic_mem_counter[288] = 4'b0000;
    GSharePlugin_logic_mem_counter[289] = 4'b0000;
    GSharePlugin_logic_mem_counter[290] = 4'b0000;
    GSharePlugin_logic_mem_counter[291] = 4'b0000;
    GSharePlugin_logic_mem_counter[292] = 4'b0000;
    GSharePlugin_logic_mem_counter[293] = 4'b0000;
    GSharePlugin_logic_mem_counter[294] = 4'b0000;
    GSharePlugin_logic_mem_counter[295] = 4'b0000;
    GSharePlugin_logic_mem_counter[296] = 4'b0000;
    GSharePlugin_logic_mem_counter[297] = 4'b0000;
    GSharePlugin_logic_mem_counter[298] = 4'b0000;
    GSharePlugin_logic_mem_counter[299] = 4'b0000;
    GSharePlugin_logic_mem_counter[300] = 4'b0000;
    GSharePlugin_logic_mem_counter[301] = 4'b0000;
    GSharePlugin_logic_mem_counter[302] = 4'b0000;
    GSharePlugin_logic_mem_counter[303] = 4'b0000;
    GSharePlugin_logic_mem_counter[304] = 4'b0000;
    GSharePlugin_logic_mem_counter[305] = 4'b0000;
    GSharePlugin_logic_mem_counter[306] = 4'b0000;
    GSharePlugin_logic_mem_counter[307] = 4'b0000;
    GSharePlugin_logic_mem_counter[308] = 4'b0000;
    GSharePlugin_logic_mem_counter[309] = 4'b0000;
    GSharePlugin_logic_mem_counter[310] = 4'b0000;
    GSharePlugin_logic_mem_counter[311] = 4'b0000;
    GSharePlugin_logic_mem_counter[312] = 4'b0000;
    GSharePlugin_logic_mem_counter[313] = 4'b0000;
    GSharePlugin_logic_mem_counter[314] = 4'b0000;
    GSharePlugin_logic_mem_counter[315] = 4'b0000;
    GSharePlugin_logic_mem_counter[316] = 4'b0000;
    GSharePlugin_logic_mem_counter[317] = 4'b0000;
    GSharePlugin_logic_mem_counter[318] = 4'b0000;
    GSharePlugin_logic_mem_counter[319] = 4'b0000;
    GSharePlugin_logic_mem_counter[320] = 4'b0000;
    GSharePlugin_logic_mem_counter[321] = 4'b0000;
    GSharePlugin_logic_mem_counter[322] = 4'b0000;
    GSharePlugin_logic_mem_counter[323] = 4'b0000;
    GSharePlugin_logic_mem_counter[324] = 4'b0000;
    GSharePlugin_logic_mem_counter[325] = 4'b0000;
    GSharePlugin_logic_mem_counter[326] = 4'b0000;
    GSharePlugin_logic_mem_counter[327] = 4'b0000;
    GSharePlugin_logic_mem_counter[328] = 4'b0000;
    GSharePlugin_logic_mem_counter[329] = 4'b0000;
    GSharePlugin_logic_mem_counter[330] = 4'b0000;
    GSharePlugin_logic_mem_counter[331] = 4'b0000;
    GSharePlugin_logic_mem_counter[332] = 4'b0000;
    GSharePlugin_logic_mem_counter[333] = 4'b0000;
    GSharePlugin_logic_mem_counter[334] = 4'b0000;
    GSharePlugin_logic_mem_counter[335] = 4'b0000;
    GSharePlugin_logic_mem_counter[336] = 4'b0000;
    GSharePlugin_logic_mem_counter[337] = 4'b0000;
    GSharePlugin_logic_mem_counter[338] = 4'b0000;
    GSharePlugin_logic_mem_counter[339] = 4'b0000;
    GSharePlugin_logic_mem_counter[340] = 4'b0000;
    GSharePlugin_logic_mem_counter[341] = 4'b0000;
    GSharePlugin_logic_mem_counter[342] = 4'b0000;
    GSharePlugin_logic_mem_counter[343] = 4'b0000;
    GSharePlugin_logic_mem_counter[344] = 4'b0000;
    GSharePlugin_logic_mem_counter[345] = 4'b0000;
    GSharePlugin_logic_mem_counter[346] = 4'b0000;
    GSharePlugin_logic_mem_counter[347] = 4'b0000;
    GSharePlugin_logic_mem_counter[348] = 4'b0000;
    GSharePlugin_logic_mem_counter[349] = 4'b0000;
    GSharePlugin_logic_mem_counter[350] = 4'b0000;
    GSharePlugin_logic_mem_counter[351] = 4'b0000;
    GSharePlugin_logic_mem_counter[352] = 4'b0000;
    GSharePlugin_logic_mem_counter[353] = 4'b0000;
    GSharePlugin_logic_mem_counter[354] = 4'b0000;
    GSharePlugin_logic_mem_counter[355] = 4'b0000;
    GSharePlugin_logic_mem_counter[356] = 4'b0000;
    GSharePlugin_logic_mem_counter[357] = 4'b0000;
    GSharePlugin_logic_mem_counter[358] = 4'b0000;
    GSharePlugin_logic_mem_counter[359] = 4'b0000;
    GSharePlugin_logic_mem_counter[360] = 4'b0000;
    GSharePlugin_logic_mem_counter[361] = 4'b0000;
    GSharePlugin_logic_mem_counter[362] = 4'b0000;
    GSharePlugin_logic_mem_counter[363] = 4'b0000;
    GSharePlugin_logic_mem_counter[364] = 4'b0000;
    GSharePlugin_logic_mem_counter[365] = 4'b0000;
    GSharePlugin_logic_mem_counter[366] = 4'b0000;
    GSharePlugin_logic_mem_counter[367] = 4'b0000;
    GSharePlugin_logic_mem_counter[368] = 4'b0000;
    GSharePlugin_logic_mem_counter[369] = 4'b0000;
    GSharePlugin_logic_mem_counter[370] = 4'b0000;
    GSharePlugin_logic_mem_counter[371] = 4'b0000;
    GSharePlugin_logic_mem_counter[372] = 4'b0000;
    GSharePlugin_logic_mem_counter[373] = 4'b0000;
    GSharePlugin_logic_mem_counter[374] = 4'b0000;
    GSharePlugin_logic_mem_counter[375] = 4'b0000;
    GSharePlugin_logic_mem_counter[376] = 4'b0000;
    GSharePlugin_logic_mem_counter[377] = 4'b0000;
    GSharePlugin_logic_mem_counter[378] = 4'b0000;
    GSharePlugin_logic_mem_counter[379] = 4'b0000;
    GSharePlugin_logic_mem_counter[380] = 4'b0000;
    GSharePlugin_logic_mem_counter[381] = 4'b0000;
    GSharePlugin_logic_mem_counter[382] = 4'b0000;
    GSharePlugin_logic_mem_counter[383] = 4'b0000;
    GSharePlugin_logic_mem_counter[384] = 4'b0000;
    GSharePlugin_logic_mem_counter[385] = 4'b0000;
    GSharePlugin_logic_mem_counter[386] = 4'b0000;
    GSharePlugin_logic_mem_counter[387] = 4'b0000;
    GSharePlugin_logic_mem_counter[388] = 4'b0000;
    GSharePlugin_logic_mem_counter[389] = 4'b0000;
    GSharePlugin_logic_mem_counter[390] = 4'b0000;
    GSharePlugin_logic_mem_counter[391] = 4'b0000;
    GSharePlugin_logic_mem_counter[392] = 4'b0000;
    GSharePlugin_logic_mem_counter[393] = 4'b0000;
    GSharePlugin_logic_mem_counter[394] = 4'b0000;
    GSharePlugin_logic_mem_counter[395] = 4'b0000;
    GSharePlugin_logic_mem_counter[396] = 4'b0000;
    GSharePlugin_logic_mem_counter[397] = 4'b0000;
    GSharePlugin_logic_mem_counter[398] = 4'b0000;
    GSharePlugin_logic_mem_counter[399] = 4'b0000;
    GSharePlugin_logic_mem_counter[400] = 4'b0000;
    GSharePlugin_logic_mem_counter[401] = 4'b0000;
    GSharePlugin_logic_mem_counter[402] = 4'b0000;
    GSharePlugin_logic_mem_counter[403] = 4'b0000;
    GSharePlugin_logic_mem_counter[404] = 4'b0000;
    GSharePlugin_logic_mem_counter[405] = 4'b0000;
    GSharePlugin_logic_mem_counter[406] = 4'b0000;
    GSharePlugin_logic_mem_counter[407] = 4'b0000;
    GSharePlugin_logic_mem_counter[408] = 4'b0000;
    GSharePlugin_logic_mem_counter[409] = 4'b0000;
    GSharePlugin_logic_mem_counter[410] = 4'b0000;
    GSharePlugin_logic_mem_counter[411] = 4'b0000;
    GSharePlugin_logic_mem_counter[412] = 4'b0000;
    GSharePlugin_logic_mem_counter[413] = 4'b0000;
    GSharePlugin_logic_mem_counter[414] = 4'b0000;
    GSharePlugin_logic_mem_counter[415] = 4'b0000;
    GSharePlugin_logic_mem_counter[416] = 4'b0000;
    GSharePlugin_logic_mem_counter[417] = 4'b0000;
    GSharePlugin_logic_mem_counter[418] = 4'b0000;
    GSharePlugin_logic_mem_counter[419] = 4'b0000;
    GSharePlugin_logic_mem_counter[420] = 4'b0000;
    GSharePlugin_logic_mem_counter[421] = 4'b0000;
    GSharePlugin_logic_mem_counter[422] = 4'b0000;
    GSharePlugin_logic_mem_counter[423] = 4'b0000;
    GSharePlugin_logic_mem_counter[424] = 4'b0000;
    GSharePlugin_logic_mem_counter[425] = 4'b0000;
    GSharePlugin_logic_mem_counter[426] = 4'b0000;
    GSharePlugin_logic_mem_counter[427] = 4'b0000;
    GSharePlugin_logic_mem_counter[428] = 4'b0000;
    GSharePlugin_logic_mem_counter[429] = 4'b0000;
    GSharePlugin_logic_mem_counter[430] = 4'b0000;
    GSharePlugin_logic_mem_counter[431] = 4'b0000;
    GSharePlugin_logic_mem_counter[432] = 4'b0000;
    GSharePlugin_logic_mem_counter[433] = 4'b0000;
    GSharePlugin_logic_mem_counter[434] = 4'b0000;
    GSharePlugin_logic_mem_counter[435] = 4'b0000;
    GSharePlugin_logic_mem_counter[436] = 4'b0000;
    GSharePlugin_logic_mem_counter[437] = 4'b0000;
    GSharePlugin_logic_mem_counter[438] = 4'b0000;
    GSharePlugin_logic_mem_counter[439] = 4'b0000;
    GSharePlugin_logic_mem_counter[440] = 4'b0000;
    GSharePlugin_logic_mem_counter[441] = 4'b0000;
    GSharePlugin_logic_mem_counter[442] = 4'b0000;
    GSharePlugin_logic_mem_counter[443] = 4'b0000;
    GSharePlugin_logic_mem_counter[444] = 4'b0000;
    GSharePlugin_logic_mem_counter[445] = 4'b0000;
    GSharePlugin_logic_mem_counter[446] = 4'b0000;
    GSharePlugin_logic_mem_counter[447] = 4'b0000;
    GSharePlugin_logic_mem_counter[448] = 4'b0000;
    GSharePlugin_logic_mem_counter[449] = 4'b0000;
    GSharePlugin_logic_mem_counter[450] = 4'b0000;
    GSharePlugin_logic_mem_counter[451] = 4'b0000;
    GSharePlugin_logic_mem_counter[452] = 4'b0000;
    GSharePlugin_logic_mem_counter[453] = 4'b0000;
    GSharePlugin_logic_mem_counter[454] = 4'b0000;
    GSharePlugin_logic_mem_counter[455] = 4'b0000;
    GSharePlugin_logic_mem_counter[456] = 4'b0000;
    GSharePlugin_logic_mem_counter[457] = 4'b0000;
    GSharePlugin_logic_mem_counter[458] = 4'b0000;
    GSharePlugin_logic_mem_counter[459] = 4'b0000;
    GSharePlugin_logic_mem_counter[460] = 4'b0000;
    GSharePlugin_logic_mem_counter[461] = 4'b0000;
    GSharePlugin_logic_mem_counter[462] = 4'b0000;
    GSharePlugin_logic_mem_counter[463] = 4'b0000;
    GSharePlugin_logic_mem_counter[464] = 4'b0000;
    GSharePlugin_logic_mem_counter[465] = 4'b0000;
    GSharePlugin_logic_mem_counter[466] = 4'b0000;
    GSharePlugin_logic_mem_counter[467] = 4'b0000;
    GSharePlugin_logic_mem_counter[468] = 4'b0000;
    GSharePlugin_logic_mem_counter[469] = 4'b0000;
    GSharePlugin_logic_mem_counter[470] = 4'b0000;
    GSharePlugin_logic_mem_counter[471] = 4'b0000;
    GSharePlugin_logic_mem_counter[472] = 4'b0000;
    GSharePlugin_logic_mem_counter[473] = 4'b0000;
    GSharePlugin_logic_mem_counter[474] = 4'b0000;
    GSharePlugin_logic_mem_counter[475] = 4'b0000;
    GSharePlugin_logic_mem_counter[476] = 4'b0000;
    GSharePlugin_logic_mem_counter[477] = 4'b0000;
    GSharePlugin_logic_mem_counter[478] = 4'b0000;
    GSharePlugin_logic_mem_counter[479] = 4'b0000;
    GSharePlugin_logic_mem_counter[480] = 4'b0000;
    GSharePlugin_logic_mem_counter[481] = 4'b0000;
    GSharePlugin_logic_mem_counter[482] = 4'b0000;
    GSharePlugin_logic_mem_counter[483] = 4'b0000;
    GSharePlugin_logic_mem_counter[484] = 4'b0000;
    GSharePlugin_logic_mem_counter[485] = 4'b0000;
    GSharePlugin_logic_mem_counter[486] = 4'b0000;
    GSharePlugin_logic_mem_counter[487] = 4'b0000;
    GSharePlugin_logic_mem_counter[488] = 4'b0000;
    GSharePlugin_logic_mem_counter[489] = 4'b0000;
    GSharePlugin_logic_mem_counter[490] = 4'b0000;
    GSharePlugin_logic_mem_counter[491] = 4'b0000;
    GSharePlugin_logic_mem_counter[492] = 4'b0000;
    GSharePlugin_logic_mem_counter[493] = 4'b0000;
    GSharePlugin_logic_mem_counter[494] = 4'b0000;
    GSharePlugin_logic_mem_counter[495] = 4'b0000;
    GSharePlugin_logic_mem_counter[496] = 4'b0000;
    GSharePlugin_logic_mem_counter[497] = 4'b0000;
    GSharePlugin_logic_mem_counter[498] = 4'b0000;
    GSharePlugin_logic_mem_counter[499] = 4'b0000;
    GSharePlugin_logic_mem_counter[500] = 4'b0000;
    GSharePlugin_logic_mem_counter[501] = 4'b0000;
    GSharePlugin_logic_mem_counter[502] = 4'b0000;
    GSharePlugin_logic_mem_counter[503] = 4'b0000;
    GSharePlugin_logic_mem_counter[504] = 4'b0000;
    GSharePlugin_logic_mem_counter[505] = 4'b0000;
    GSharePlugin_logic_mem_counter[506] = 4'b0000;
    GSharePlugin_logic_mem_counter[507] = 4'b0000;
    GSharePlugin_logic_mem_counter[508] = 4'b0000;
    GSharePlugin_logic_mem_counter[509] = 4'b0000;
    GSharePlugin_logic_mem_counter[510] = 4'b0000;
    GSharePlugin_logic_mem_counter[511] = 4'b0000;
    GSharePlugin_logic_mem_counter[512] = 4'b0000;
    GSharePlugin_logic_mem_counter[513] = 4'b0000;
    GSharePlugin_logic_mem_counter[514] = 4'b0000;
    GSharePlugin_logic_mem_counter[515] = 4'b0000;
    GSharePlugin_logic_mem_counter[516] = 4'b0000;
    GSharePlugin_logic_mem_counter[517] = 4'b0000;
    GSharePlugin_logic_mem_counter[518] = 4'b0000;
    GSharePlugin_logic_mem_counter[519] = 4'b0000;
    GSharePlugin_logic_mem_counter[520] = 4'b0000;
    GSharePlugin_logic_mem_counter[521] = 4'b0000;
    GSharePlugin_logic_mem_counter[522] = 4'b0000;
    GSharePlugin_logic_mem_counter[523] = 4'b0000;
    GSharePlugin_logic_mem_counter[524] = 4'b0000;
    GSharePlugin_logic_mem_counter[525] = 4'b0000;
    GSharePlugin_logic_mem_counter[526] = 4'b0000;
    GSharePlugin_logic_mem_counter[527] = 4'b0000;
    GSharePlugin_logic_mem_counter[528] = 4'b0000;
    GSharePlugin_logic_mem_counter[529] = 4'b0000;
    GSharePlugin_logic_mem_counter[530] = 4'b0000;
    GSharePlugin_logic_mem_counter[531] = 4'b0000;
    GSharePlugin_logic_mem_counter[532] = 4'b0000;
    GSharePlugin_logic_mem_counter[533] = 4'b0000;
    GSharePlugin_logic_mem_counter[534] = 4'b0000;
    GSharePlugin_logic_mem_counter[535] = 4'b0000;
    GSharePlugin_logic_mem_counter[536] = 4'b0000;
    GSharePlugin_logic_mem_counter[537] = 4'b0000;
    GSharePlugin_logic_mem_counter[538] = 4'b0000;
    GSharePlugin_logic_mem_counter[539] = 4'b0000;
    GSharePlugin_logic_mem_counter[540] = 4'b0000;
    GSharePlugin_logic_mem_counter[541] = 4'b0000;
    GSharePlugin_logic_mem_counter[542] = 4'b0000;
    GSharePlugin_logic_mem_counter[543] = 4'b0000;
    GSharePlugin_logic_mem_counter[544] = 4'b0000;
    GSharePlugin_logic_mem_counter[545] = 4'b0000;
    GSharePlugin_logic_mem_counter[546] = 4'b0000;
    GSharePlugin_logic_mem_counter[547] = 4'b0000;
    GSharePlugin_logic_mem_counter[548] = 4'b0000;
    GSharePlugin_logic_mem_counter[549] = 4'b0000;
    GSharePlugin_logic_mem_counter[550] = 4'b0000;
    GSharePlugin_logic_mem_counter[551] = 4'b0000;
    GSharePlugin_logic_mem_counter[552] = 4'b0000;
    GSharePlugin_logic_mem_counter[553] = 4'b0000;
    GSharePlugin_logic_mem_counter[554] = 4'b0000;
    GSharePlugin_logic_mem_counter[555] = 4'b0000;
    GSharePlugin_logic_mem_counter[556] = 4'b0000;
    GSharePlugin_logic_mem_counter[557] = 4'b0000;
    GSharePlugin_logic_mem_counter[558] = 4'b0000;
    GSharePlugin_logic_mem_counter[559] = 4'b0000;
    GSharePlugin_logic_mem_counter[560] = 4'b0000;
    GSharePlugin_logic_mem_counter[561] = 4'b0000;
    GSharePlugin_logic_mem_counter[562] = 4'b0000;
    GSharePlugin_logic_mem_counter[563] = 4'b0000;
    GSharePlugin_logic_mem_counter[564] = 4'b0000;
    GSharePlugin_logic_mem_counter[565] = 4'b0000;
    GSharePlugin_logic_mem_counter[566] = 4'b0000;
    GSharePlugin_logic_mem_counter[567] = 4'b0000;
    GSharePlugin_logic_mem_counter[568] = 4'b0000;
    GSharePlugin_logic_mem_counter[569] = 4'b0000;
    GSharePlugin_logic_mem_counter[570] = 4'b0000;
    GSharePlugin_logic_mem_counter[571] = 4'b0000;
    GSharePlugin_logic_mem_counter[572] = 4'b0000;
    GSharePlugin_logic_mem_counter[573] = 4'b0000;
    GSharePlugin_logic_mem_counter[574] = 4'b0000;
    GSharePlugin_logic_mem_counter[575] = 4'b0000;
    GSharePlugin_logic_mem_counter[576] = 4'b0000;
    GSharePlugin_logic_mem_counter[577] = 4'b0000;
    GSharePlugin_logic_mem_counter[578] = 4'b0000;
    GSharePlugin_logic_mem_counter[579] = 4'b0000;
    GSharePlugin_logic_mem_counter[580] = 4'b0000;
    GSharePlugin_logic_mem_counter[581] = 4'b0000;
    GSharePlugin_logic_mem_counter[582] = 4'b0000;
    GSharePlugin_logic_mem_counter[583] = 4'b0000;
    GSharePlugin_logic_mem_counter[584] = 4'b0000;
    GSharePlugin_logic_mem_counter[585] = 4'b0000;
    GSharePlugin_logic_mem_counter[586] = 4'b0000;
    GSharePlugin_logic_mem_counter[587] = 4'b0000;
    GSharePlugin_logic_mem_counter[588] = 4'b0000;
    GSharePlugin_logic_mem_counter[589] = 4'b0000;
    GSharePlugin_logic_mem_counter[590] = 4'b0000;
    GSharePlugin_logic_mem_counter[591] = 4'b0000;
    GSharePlugin_logic_mem_counter[592] = 4'b0000;
    GSharePlugin_logic_mem_counter[593] = 4'b0000;
    GSharePlugin_logic_mem_counter[594] = 4'b0000;
    GSharePlugin_logic_mem_counter[595] = 4'b0000;
    GSharePlugin_logic_mem_counter[596] = 4'b0000;
    GSharePlugin_logic_mem_counter[597] = 4'b0000;
    GSharePlugin_logic_mem_counter[598] = 4'b0000;
    GSharePlugin_logic_mem_counter[599] = 4'b0000;
    GSharePlugin_logic_mem_counter[600] = 4'b0000;
    GSharePlugin_logic_mem_counter[601] = 4'b0000;
    GSharePlugin_logic_mem_counter[602] = 4'b0000;
    GSharePlugin_logic_mem_counter[603] = 4'b0000;
    GSharePlugin_logic_mem_counter[604] = 4'b0000;
    GSharePlugin_logic_mem_counter[605] = 4'b0000;
    GSharePlugin_logic_mem_counter[606] = 4'b0000;
    GSharePlugin_logic_mem_counter[607] = 4'b0000;
    GSharePlugin_logic_mem_counter[608] = 4'b0000;
    GSharePlugin_logic_mem_counter[609] = 4'b0000;
    GSharePlugin_logic_mem_counter[610] = 4'b0000;
    GSharePlugin_logic_mem_counter[611] = 4'b0000;
    GSharePlugin_logic_mem_counter[612] = 4'b0000;
    GSharePlugin_logic_mem_counter[613] = 4'b0000;
    GSharePlugin_logic_mem_counter[614] = 4'b0000;
    GSharePlugin_logic_mem_counter[615] = 4'b0000;
    GSharePlugin_logic_mem_counter[616] = 4'b0000;
    GSharePlugin_logic_mem_counter[617] = 4'b0000;
    GSharePlugin_logic_mem_counter[618] = 4'b0000;
    GSharePlugin_logic_mem_counter[619] = 4'b0000;
    GSharePlugin_logic_mem_counter[620] = 4'b0000;
    GSharePlugin_logic_mem_counter[621] = 4'b0000;
    GSharePlugin_logic_mem_counter[622] = 4'b0000;
    GSharePlugin_logic_mem_counter[623] = 4'b0000;
    GSharePlugin_logic_mem_counter[624] = 4'b0000;
    GSharePlugin_logic_mem_counter[625] = 4'b0000;
    GSharePlugin_logic_mem_counter[626] = 4'b0000;
    GSharePlugin_logic_mem_counter[627] = 4'b0000;
    GSharePlugin_logic_mem_counter[628] = 4'b0000;
    GSharePlugin_logic_mem_counter[629] = 4'b0000;
    GSharePlugin_logic_mem_counter[630] = 4'b0000;
    GSharePlugin_logic_mem_counter[631] = 4'b0000;
    GSharePlugin_logic_mem_counter[632] = 4'b0000;
    GSharePlugin_logic_mem_counter[633] = 4'b0000;
    GSharePlugin_logic_mem_counter[634] = 4'b0000;
    GSharePlugin_logic_mem_counter[635] = 4'b0000;
    GSharePlugin_logic_mem_counter[636] = 4'b0000;
    GSharePlugin_logic_mem_counter[637] = 4'b0000;
    GSharePlugin_logic_mem_counter[638] = 4'b0000;
    GSharePlugin_logic_mem_counter[639] = 4'b0000;
    GSharePlugin_logic_mem_counter[640] = 4'b0000;
    GSharePlugin_logic_mem_counter[641] = 4'b0000;
    GSharePlugin_logic_mem_counter[642] = 4'b0000;
    GSharePlugin_logic_mem_counter[643] = 4'b0000;
    GSharePlugin_logic_mem_counter[644] = 4'b0000;
    GSharePlugin_logic_mem_counter[645] = 4'b0000;
    GSharePlugin_logic_mem_counter[646] = 4'b0000;
    GSharePlugin_logic_mem_counter[647] = 4'b0000;
    GSharePlugin_logic_mem_counter[648] = 4'b0000;
    GSharePlugin_logic_mem_counter[649] = 4'b0000;
    GSharePlugin_logic_mem_counter[650] = 4'b0000;
    GSharePlugin_logic_mem_counter[651] = 4'b0000;
    GSharePlugin_logic_mem_counter[652] = 4'b0000;
    GSharePlugin_logic_mem_counter[653] = 4'b0000;
    GSharePlugin_logic_mem_counter[654] = 4'b0000;
    GSharePlugin_logic_mem_counter[655] = 4'b0000;
    GSharePlugin_logic_mem_counter[656] = 4'b0000;
    GSharePlugin_logic_mem_counter[657] = 4'b0000;
    GSharePlugin_logic_mem_counter[658] = 4'b0000;
    GSharePlugin_logic_mem_counter[659] = 4'b0000;
    GSharePlugin_logic_mem_counter[660] = 4'b0000;
    GSharePlugin_logic_mem_counter[661] = 4'b0000;
    GSharePlugin_logic_mem_counter[662] = 4'b0000;
    GSharePlugin_logic_mem_counter[663] = 4'b0000;
    GSharePlugin_logic_mem_counter[664] = 4'b0000;
    GSharePlugin_logic_mem_counter[665] = 4'b0000;
    GSharePlugin_logic_mem_counter[666] = 4'b0000;
    GSharePlugin_logic_mem_counter[667] = 4'b0000;
    GSharePlugin_logic_mem_counter[668] = 4'b0000;
    GSharePlugin_logic_mem_counter[669] = 4'b0000;
    GSharePlugin_logic_mem_counter[670] = 4'b0000;
    GSharePlugin_logic_mem_counter[671] = 4'b0000;
    GSharePlugin_logic_mem_counter[672] = 4'b0000;
    GSharePlugin_logic_mem_counter[673] = 4'b0000;
    GSharePlugin_logic_mem_counter[674] = 4'b0000;
    GSharePlugin_logic_mem_counter[675] = 4'b0000;
    GSharePlugin_logic_mem_counter[676] = 4'b0000;
    GSharePlugin_logic_mem_counter[677] = 4'b0000;
    GSharePlugin_logic_mem_counter[678] = 4'b0000;
    GSharePlugin_logic_mem_counter[679] = 4'b0000;
    GSharePlugin_logic_mem_counter[680] = 4'b0000;
    GSharePlugin_logic_mem_counter[681] = 4'b0000;
    GSharePlugin_logic_mem_counter[682] = 4'b0000;
    GSharePlugin_logic_mem_counter[683] = 4'b0000;
    GSharePlugin_logic_mem_counter[684] = 4'b0000;
    GSharePlugin_logic_mem_counter[685] = 4'b0000;
    GSharePlugin_logic_mem_counter[686] = 4'b0000;
    GSharePlugin_logic_mem_counter[687] = 4'b0000;
    GSharePlugin_logic_mem_counter[688] = 4'b0000;
    GSharePlugin_logic_mem_counter[689] = 4'b0000;
    GSharePlugin_logic_mem_counter[690] = 4'b0000;
    GSharePlugin_logic_mem_counter[691] = 4'b0000;
    GSharePlugin_logic_mem_counter[692] = 4'b0000;
    GSharePlugin_logic_mem_counter[693] = 4'b0000;
    GSharePlugin_logic_mem_counter[694] = 4'b0000;
    GSharePlugin_logic_mem_counter[695] = 4'b0000;
    GSharePlugin_logic_mem_counter[696] = 4'b0000;
    GSharePlugin_logic_mem_counter[697] = 4'b0000;
    GSharePlugin_logic_mem_counter[698] = 4'b0000;
    GSharePlugin_logic_mem_counter[699] = 4'b0000;
    GSharePlugin_logic_mem_counter[700] = 4'b0000;
    GSharePlugin_logic_mem_counter[701] = 4'b0000;
    GSharePlugin_logic_mem_counter[702] = 4'b0000;
    GSharePlugin_logic_mem_counter[703] = 4'b0000;
    GSharePlugin_logic_mem_counter[704] = 4'b0000;
    GSharePlugin_logic_mem_counter[705] = 4'b0000;
    GSharePlugin_logic_mem_counter[706] = 4'b0000;
    GSharePlugin_logic_mem_counter[707] = 4'b0000;
    GSharePlugin_logic_mem_counter[708] = 4'b0000;
    GSharePlugin_logic_mem_counter[709] = 4'b0000;
    GSharePlugin_logic_mem_counter[710] = 4'b0000;
    GSharePlugin_logic_mem_counter[711] = 4'b0000;
    GSharePlugin_logic_mem_counter[712] = 4'b0000;
    GSharePlugin_logic_mem_counter[713] = 4'b0000;
    GSharePlugin_logic_mem_counter[714] = 4'b0000;
    GSharePlugin_logic_mem_counter[715] = 4'b0000;
    GSharePlugin_logic_mem_counter[716] = 4'b0000;
    GSharePlugin_logic_mem_counter[717] = 4'b0000;
    GSharePlugin_logic_mem_counter[718] = 4'b0000;
    GSharePlugin_logic_mem_counter[719] = 4'b0000;
    GSharePlugin_logic_mem_counter[720] = 4'b0000;
    GSharePlugin_logic_mem_counter[721] = 4'b0000;
    GSharePlugin_logic_mem_counter[722] = 4'b0000;
    GSharePlugin_logic_mem_counter[723] = 4'b0000;
    GSharePlugin_logic_mem_counter[724] = 4'b0000;
    GSharePlugin_logic_mem_counter[725] = 4'b0000;
    GSharePlugin_logic_mem_counter[726] = 4'b0000;
    GSharePlugin_logic_mem_counter[727] = 4'b0000;
    GSharePlugin_logic_mem_counter[728] = 4'b0000;
    GSharePlugin_logic_mem_counter[729] = 4'b0000;
    GSharePlugin_logic_mem_counter[730] = 4'b0000;
    GSharePlugin_logic_mem_counter[731] = 4'b0000;
    GSharePlugin_logic_mem_counter[732] = 4'b0000;
    GSharePlugin_logic_mem_counter[733] = 4'b0000;
    GSharePlugin_logic_mem_counter[734] = 4'b0000;
    GSharePlugin_logic_mem_counter[735] = 4'b0000;
    GSharePlugin_logic_mem_counter[736] = 4'b0000;
    GSharePlugin_logic_mem_counter[737] = 4'b0000;
    GSharePlugin_logic_mem_counter[738] = 4'b0000;
    GSharePlugin_logic_mem_counter[739] = 4'b0000;
    GSharePlugin_logic_mem_counter[740] = 4'b0000;
    GSharePlugin_logic_mem_counter[741] = 4'b0000;
    GSharePlugin_logic_mem_counter[742] = 4'b0000;
    GSharePlugin_logic_mem_counter[743] = 4'b0000;
    GSharePlugin_logic_mem_counter[744] = 4'b0000;
    GSharePlugin_logic_mem_counter[745] = 4'b0000;
    GSharePlugin_logic_mem_counter[746] = 4'b0000;
    GSharePlugin_logic_mem_counter[747] = 4'b0000;
    GSharePlugin_logic_mem_counter[748] = 4'b0000;
    GSharePlugin_logic_mem_counter[749] = 4'b0000;
    GSharePlugin_logic_mem_counter[750] = 4'b0000;
    GSharePlugin_logic_mem_counter[751] = 4'b0000;
    GSharePlugin_logic_mem_counter[752] = 4'b0000;
    GSharePlugin_logic_mem_counter[753] = 4'b0000;
    GSharePlugin_logic_mem_counter[754] = 4'b0000;
    GSharePlugin_logic_mem_counter[755] = 4'b0000;
    GSharePlugin_logic_mem_counter[756] = 4'b0000;
    GSharePlugin_logic_mem_counter[757] = 4'b0000;
    GSharePlugin_logic_mem_counter[758] = 4'b0000;
    GSharePlugin_logic_mem_counter[759] = 4'b0000;
    GSharePlugin_logic_mem_counter[760] = 4'b0000;
    GSharePlugin_logic_mem_counter[761] = 4'b0000;
    GSharePlugin_logic_mem_counter[762] = 4'b0000;
    GSharePlugin_logic_mem_counter[763] = 4'b0000;
    GSharePlugin_logic_mem_counter[764] = 4'b0000;
    GSharePlugin_logic_mem_counter[765] = 4'b0000;
    GSharePlugin_logic_mem_counter[766] = 4'b0000;
    GSharePlugin_logic_mem_counter[767] = 4'b0000;
    GSharePlugin_logic_mem_counter[768] = 4'b0000;
    GSharePlugin_logic_mem_counter[769] = 4'b0000;
    GSharePlugin_logic_mem_counter[770] = 4'b0000;
    GSharePlugin_logic_mem_counter[771] = 4'b0000;
    GSharePlugin_logic_mem_counter[772] = 4'b0000;
    GSharePlugin_logic_mem_counter[773] = 4'b0000;
    GSharePlugin_logic_mem_counter[774] = 4'b0000;
    GSharePlugin_logic_mem_counter[775] = 4'b0000;
    GSharePlugin_logic_mem_counter[776] = 4'b0000;
    GSharePlugin_logic_mem_counter[777] = 4'b0000;
    GSharePlugin_logic_mem_counter[778] = 4'b0000;
    GSharePlugin_logic_mem_counter[779] = 4'b0000;
    GSharePlugin_logic_mem_counter[780] = 4'b0000;
    GSharePlugin_logic_mem_counter[781] = 4'b0000;
    GSharePlugin_logic_mem_counter[782] = 4'b0000;
    GSharePlugin_logic_mem_counter[783] = 4'b0000;
    GSharePlugin_logic_mem_counter[784] = 4'b0000;
    GSharePlugin_logic_mem_counter[785] = 4'b0000;
    GSharePlugin_logic_mem_counter[786] = 4'b0000;
    GSharePlugin_logic_mem_counter[787] = 4'b0000;
    GSharePlugin_logic_mem_counter[788] = 4'b0000;
    GSharePlugin_logic_mem_counter[789] = 4'b0000;
    GSharePlugin_logic_mem_counter[790] = 4'b0000;
    GSharePlugin_logic_mem_counter[791] = 4'b0000;
    GSharePlugin_logic_mem_counter[792] = 4'b0000;
    GSharePlugin_logic_mem_counter[793] = 4'b0000;
    GSharePlugin_logic_mem_counter[794] = 4'b0000;
    GSharePlugin_logic_mem_counter[795] = 4'b0000;
    GSharePlugin_logic_mem_counter[796] = 4'b0000;
    GSharePlugin_logic_mem_counter[797] = 4'b0000;
    GSharePlugin_logic_mem_counter[798] = 4'b0000;
    GSharePlugin_logic_mem_counter[799] = 4'b0000;
    GSharePlugin_logic_mem_counter[800] = 4'b0000;
    GSharePlugin_logic_mem_counter[801] = 4'b0000;
    GSharePlugin_logic_mem_counter[802] = 4'b0000;
    GSharePlugin_logic_mem_counter[803] = 4'b0000;
    GSharePlugin_logic_mem_counter[804] = 4'b0000;
    GSharePlugin_logic_mem_counter[805] = 4'b0000;
    GSharePlugin_logic_mem_counter[806] = 4'b0000;
    GSharePlugin_logic_mem_counter[807] = 4'b0000;
    GSharePlugin_logic_mem_counter[808] = 4'b0000;
    GSharePlugin_logic_mem_counter[809] = 4'b0000;
    GSharePlugin_logic_mem_counter[810] = 4'b0000;
    GSharePlugin_logic_mem_counter[811] = 4'b0000;
    GSharePlugin_logic_mem_counter[812] = 4'b0000;
    GSharePlugin_logic_mem_counter[813] = 4'b0000;
    GSharePlugin_logic_mem_counter[814] = 4'b0000;
    GSharePlugin_logic_mem_counter[815] = 4'b0000;
    GSharePlugin_logic_mem_counter[816] = 4'b0000;
    GSharePlugin_logic_mem_counter[817] = 4'b0000;
    GSharePlugin_logic_mem_counter[818] = 4'b0000;
    GSharePlugin_logic_mem_counter[819] = 4'b0000;
    GSharePlugin_logic_mem_counter[820] = 4'b0000;
    GSharePlugin_logic_mem_counter[821] = 4'b0000;
    GSharePlugin_logic_mem_counter[822] = 4'b0000;
    GSharePlugin_logic_mem_counter[823] = 4'b0000;
    GSharePlugin_logic_mem_counter[824] = 4'b0000;
    GSharePlugin_logic_mem_counter[825] = 4'b0000;
    GSharePlugin_logic_mem_counter[826] = 4'b0000;
    GSharePlugin_logic_mem_counter[827] = 4'b0000;
    GSharePlugin_logic_mem_counter[828] = 4'b0000;
    GSharePlugin_logic_mem_counter[829] = 4'b0000;
    GSharePlugin_logic_mem_counter[830] = 4'b0000;
    GSharePlugin_logic_mem_counter[831] = 4'b0000;
    GSharePlugin_logic_mem_counter[832] = 4'b0000;
    GSharePlugin_logic_mem_counter[833] = 4'b0000;
    GSharePlugin_logic_mem_counter[834] = 4'b0000;
    GSharePlugin_logic_mem_counter[835] = 4'b0000;
    GSharePlugin_logic_mem_counter[836] = 4'b0000;
    GSharePlugin_logic_mem_counter[837] = 4'b0000;
    GSharePlugin_logic_mem_counter[838] = 4'b0000;
    GSharePlugin_logic_mem_counter[839] = 4'b0000;
    GSharePlugin_logic_mem_counter[840] = 4'b0000;
    GSharePlugin_logic_mem_counter[841] = 4'b0000;
    GSharePlugin_logic_mem_counter[842] = 4'b0000;
    GSharePlugin_logic_mem_counter[843] = 4'b0000;
    GSharePlugin_logic_mem_counter[844] = 4'b0000;
    GSharePlugin_logic_mem_counter[845] = 4'b0000;
    GSharePlugin_logic_mem_counter[846] = 4'b0000;
    GSharePlugin_logic_mem_counter[847] = 4'b0000;
    GSharePlugin_logic_mem_counter[848] = 4'b0000;
    GSharePlugin_logic_mem_counter[849] = 4'b0000;
    GSharePlugin_logic_mem_counter[850] = 4'b0000;
    GSharePlugin_logic_mem_counter[851] = 4'b0000;
    GSharePlugin_logic_mem_counter[852] = 4'b0000;
    GSharePlugin_logic_mem_counter[853] = 4'b0000;
    GSharePlugin_logic_mem_counter[854] = 4'b0000;
    GSharePlugin_logic_mem_counter[855] = 4'b0000;
    GSharePlugin_logic_mem_counter[856] = 4'b0000;
    GSharePlugin_logic_mem_counter[857] = 4'b0000;
    GSharePlugin_logic_mem_counter[858] = 4'b0000;
    GSharePlugin_logic_mem_counter[859] = 4'b0000;
    GSharePlugin_logic_mem_counter[860] = 4'b0000;
    GSharePlugin_logic_mem_counter[861] = 4'b0000;
    GSharePlugin_logic_mem_counter[862] = 4'b0000;
    GSharePlugin_logic_mem_counter[863] = 4'b0000;
    GSharePlugin_logic_mem_counter[864] = 4'b0000;
    GSharePlugin_logic_mem_counter[865] = 4'b0000;
    GSharePlugin_logic_mem_counter[866] = 4'b0000;
    GSharePlugin_logic_mem_counter[867] = 4'b0000;
    GSharePlugin_logic_mem_counter[868] = 4'b0000;
    GSharePlugin_logic_mem_counter[869] = 4'b0000;
    GSharePlugin_logic_mem_counter[870] = 4'b0000;
    GSharePlugin_logic_mem_counter[871] = 4'b0000;
    GSharePlugin_logic_mem_counter[872] = 4'b0000;
    GSharePlugin_logic_mem_counter[873] = 4'b0000;
    GSharePlugin_logic_mem_counter[874] = 4'b0000;
    GSharePlugin_logic_mem_counter[875] = 4'b0000;
    GSharePlugin_logic_mem_counter[876] = 4'b0000;
    GSharePlugin_logic_mem_counter[877] = 4'b0000;
    GSharePlugin_logic_mem_counter[878] = 4'b0000;
    GSharePlugin_logic_mem_counter[879] = 4'b0000;
    GSharePlugin_logic_mem_counter[880] = 4'b0000;
    GSharePlugin_logic_mem_counter[881] = 4'b0000;
    GSharePlugin_logic_mem_counter[882] = 4'b0000;
    GSharePlugin_logic_mem_counter[883] = 4'b0000;
    GSharePlugin_logic_mem_counter[884] = 4'b0000;
    GSharePlugin_logic_mem_counter[885] = 4'b0000;
    GSharePlugin_logic_mem_counter[886] = 4'b0000;
    GSharePlugin_logic_mem_counter[887] = 4'b0000;
    GSharePlugin_logic_mem_counter[888] = 4'b0000;
    GSharePlugin_logic_mem_counter[889] = 4'b0000;
    GSharePlugin_logic_mem_counter[890] = 4'b0000;
    GSharePlugin_logic_mem_counter[891] = 4'b0000;
    GSharePlugin_logic_mem_counter[892] = 4'b0000;
    GSharePlugin_logic_mem_counter[893] = 4'b0000;
    GSharePlugin_logic_mem_counter[894] = 4'b0000;
    GSharePlugin_logic_mem_counter[895] = 4'b0000;
    GSharePlugin_logic_mem_counter[896] = 4'b0000;
    GSharePlugin_logic_mem_counter[897] = 4'b0000;
    GSharePlugin_logic_mem_counter[898] = 4'b0000;
    GSharePlugin_logic_mem_counter[899] = 4'b0000;
    GSharePlugin_logic_mem_counter[900] = 4'b0000;
    GSharePlugin_logic_mem_counter[901] = 4'b0000;
    GSharePlugin_logic_mem_counter[902] = 4'b0000;
    GSharePlugin_logic_mem_counter[903] = 4'b0000;
    GSharePlugin_logic_mem_counter[904] = 4'b0000;
    GSharePlugin_logic_mem_counter[905] = 4'b0000;
    GSharePlugin_logic_mem_counter[906] = 4'b0000;
    GSharePlugin_logic_mem_counter[907] = 4'b0000;
    GSharePlugin_logic_mem_counter[908] = 4'b0000;
    GSharePlugin_logic_mem_counter[909] = 4'b0000;
    GSharePlugin_logic_mem_counter[910] = 4'b0000;
    GSharePlugin_logic_mem_counter[911] = 4'b0000;
    GSharePlugin_logic_mem_counter[912] = 4'b0000;
    GSharePlugin_logic_mem_counter[913] = 4'b0000;
    GSharePlugin_logic_mem_counter[914] = 4'b0000;
    GSharePlugin_logic_mem_counter[915] = 4'b0000;
    GSharePlugin_logic_mem_counter[916] = 4'b0000;
    GSharePlugin_logic_mem_counter[917] = 4'b0000;
    GSharePlugin_logic_mem_counter[918] = 4'b0000;
    GSharePlugin_logic_mem_counter[919] = 4'b0000;
    GSharePlugin_logic_mem_counter[920] = 4'b0000;
    GSharePlugin_logic_mem_counter[921] = 4'b0000;
    GSharePlugin_logic_mem_counter[922] = 4'b0000;
    GSharePlugin_logic_mem_counter[923] = 4'b0000;
    GSharePlugin_logic_mem_counter[924] = 4'b0000;
    GSharePlugin_logic_mem_counter[925] = 4'b0000;
    GSharePlugin_logic_mem_counter[926] = 4'b0000;
    GSharePlugin_logic_mem_counter[927] = 4'b0000;
    GSharePlugin_logic_mem_counter[928] = 4'b0000;
    GSharePlugin_logic_mem_counter[929] = 4'b0000;
    GSharePlugin_logic_mem_counter[930] = 4'b0000;
    GSharePlugin_logic_mem_counter[931] = 4'b0000;
    GSharePlugin_logic_mem_counter[932] = 4'b0000;
    GSharePlugin_logic_mem_counter[933] = 4'b0000;
    GSharePlugin_logic_mem_counter[934] = 4'b0000;
    GSharePlugin_logic_mem_counter[935] = 4'b0000;
    GSharePlugin_logic_mem_counter[936] = 4'b0000;
    GSharePlugin_logic_mem_counter[937] = 4'b0000;
    GSharePlugin_logic_mem_counter[938] = 4'b0000;
    GSharePlugin_logic_mem_counter[939] = 4'b0000;
    GSharePlugin_logic_mem_counter[940] = 4'b0000;
    GSharePlugin_logic_mem_counter[941] = 4'b0000;
    GSharePlugin_logic_mem_counter[942] = 4'b0000;
    GSharePlugin_logic_mem_counter[943] = 4'b0000;
    GSharePlugin_logic_mem_counter[944] = 4'b0000;
    GSharePlugin_logic_mem_counter[945] = 4'b0000;
    GSharePlugin_logic_mem_counter[946] = 4'b0000;
    GSharePlugin_logic_mem_counter[947] = 4'b0000;
    GSharePlugin_logic_mem_counter[948] = 4'b0000;
    GSharePlugin_logic_mem_counter[949] = 4'b0000;
    GSharePlugin_logic_mem_counter[950] = 4'b0000;
    GSharePlugin_logic_mem_counter[951] = 4'b0000;
    GSharePlugin_logic_mem_counter[952] = 4'b0000;
    GSharePlugin_logic_mem_counter[953] = 4'b0000;
    GSharePlugin_logic_mem_counter[954] = 4'b0000;
    GSharePlugin_logic_mem_counter[955] = 4'b0000;
    GSharePlugin_logic_mem_counter[956] = 4'b0000;
    GSharePlugin_logic_mem_counter[957] = 4'b0000;
    GSharePlugin_logic_mem_counter[958] = 4'b0000;
    GSharePlugin_logic_mem_counter[959] = 4'b0000;
    GSharePlugin_logic_mem_counter[960] = 4'b0000;
    GSharePlugin_logic_mem_counter[961] = 4'b0000;
    GSharePlugin_logic_mem_counter[962] = 4'b0000;
    GSharePlugin_logic_mem_counter[963] = 4'b0000;
    GSharePlugin_logic_mem_counter[964] = 4'b0000;
    GSharePlugin_logic_mem_counter[965] = 4'b0000;
    GSharePlugin_logic_mem_counter[966] = 4'b0000;
    GSharePlugin_logic_mem_counter[967] = 4'b0000;
    GSharePlugin_logic_mem_counter[968] = 4'b0000;
    GSharePlugin_logic_mem_counter[969] = 4'b0000;
    GSharePlugin_logic_mem_counter[970] = 4'b0000;
    GSharePlugin_logic_mem_counter[971] = 4'b0000;
    GSharePlugin_logic_mem_counter[972] = 4'b0000;
    GSharePlugin_logic_mem_counter[973] = 4'b0000;
    GSharePlugin_logic_mem_counter[974] = 4'b0000;
    GSharePlugin_logic_mem_counter[975] = 4'b0000;
    GSharePlugin_logic_mem_counter[976] = 4'b0000;
    GSharePlugin_logic_mem_counter[977] = 4'b0000;
    GSharePlugin_logic_mem_counter[978] = 4'b0000;
    GSharePlugin_logic_mem_counter[979] = 4'b0000;
    GSharePlugin_logic_mem_counter[980] = 4'b0000;
    GSharePlugin_logic_mem_counter[981] = 4'b0000;
    GSharePlugin_logic_mem_counter[982] = 4'b0000;
    GSharePlugin_logic_mem_counter[983] = 4'b0000;
    GSharePlugin_logic_mem_counter[984] = 4'b0000;
    GSharePlugin_logic_mem_counter[985] = 4'b0000;
    GSharePlugin_logic_mem_counter[986] = 4'b0000;
    GSharePlugin_logic_mem_counter[987] = 4'b0000;
    GSharePlugin_logic_mem_counter[988] = 4'b0000;
    GSharePlugin_logic_mem_counter[989] = 4'b0000;
    GSharePlugin_logic_mem_counter[990] = 4'b0000;
    GSharePlugin_logic_mem_counter[991] = 4'b0000;
    GSharePlugin_logic_mem_counter[992] = 4'b0000;
    GSharePlugin_logic_mem_counter[993] = 4'b0000;
    GSharePlugin_logic_mem_counter[994] = 4'b0000;
    GSharePlugin_logic_mem_counter[995] = 4'b0000;
    GSharePlugin_logic_mem_counter[996] = 4'b0000;
    GSharePlugin_logic_mem_counter[997] = 4'b0000;
    GSharePlugin_logic_mem_counter[998] = 4'b0000;
    GSharePlugin_logic_mem_counter[999] = 4'b0000;
    GSharePlugin_logic_mem_counter[1000] = 4'b0000;
    GSharePlugin_logic_mem_counter[1001] = 4'b0000;
    GSharePlugin_logic_mem_counter[1002] = 4'b0000;
    GSharePlugin_logic_mem_counter[1003] = 4'b0000;
    GSharePlugin_logic_mem_counter[1004] = 4'b0000;
    GSharePlugin_logic_mem_counter[1005] = 4'b0000;
    GSharePlugin_logic_mem_counter[1006] = 4'b0000;
    GSharePlugin_logic_mem_counter[1007] = 4'b0000;
    GSharePlugin_logic_mem_counter[1008] = 4'b0000;
    GSharePlugin_logic_mem_counter[1009] = 4'b0000;
    GSharePlugin_logic_mem_counter[1010] = 4'b0000;
    GSharePlugin_logic_mem_counter[1011] = 4'b0000;
    GSharePlugin_logic_mem_counter[1012] = 4'b0000;
    GSharePlugin_logic_mem_counter[1013] = 4'b0000;
    GSharePlugin_logic_mem_counter[1014] = 4'b0000;
    GSharePlugin_logic_mem_counter[1015] = 4'b0000;
    GSharePlugin_logic_mem_counter[1016] = 4'b0000;
    GSharePlugin_logic_mem_counter[1017] = 4'b0000;
    GSharePlugin_logic_mem_counter[1018] = 4'b0000;
    GSharePlugin_logic_mem_counter[1019] = 4'b0000;
    GSharePlugin_logic_mem_counter[1020] = 4'b0000;
    GSharePlugin_logic_mem_counter[1021] = 4'b0000;
    GSharePlugin_logic_mem_counter[1022] = 4'b0000;
    GSharePlugin_logic_mem_counter[1023] = 4'b0000;
    GSharePlugin_logic_mem_counter[1024] = 4'b0000;
    GSharePlugin_logic_mem_counter[1025] = 4'b0000;
    GSharePlugin_logic_mem_counter[1026] = 4'b0000;
    GSharePlugin_logic_mem_counter[1027] = 4'b0000;
    GSharePlugin_logic_mem_counter[1028] = 4'b0000;
    GSharePlugin_logic_mem_counter[1029] = 4'b0000;
    GSharePlugin_logic_mem_counter[1030] = 4'b0000;
    GSharePlugin_logic_mem_counter[1031] = 4'b0000;
    GSharePlugin_logic_mem_counter[1032] = 4'b0000;
    GSharePlugin_logic_mem_counter[1033] = 4'b0000;
    GSharePlugin_logic_mem_counter[1034] = 4'b0000;
    GSharePlugin_logic_mem_counter[1035] = 4'b0000;
    GSharePlugin_logic_mem_counter[1036] = 4'b0000;
    GSharePlugin_logic_mem_counter[1037] = 4'b0000;
    GSharePlugin_logic_mem_counter[1038] = 4'b0000;
    GSharePlugin_logic_mem_counter[1039] = 4'b0000;
    GSharePlugin_logic_mem_counter[1040] = 4'b0000;
    GSharePlugin_logic_mem_counter[1041] = 4'b0000;
    GSharePlugin_logic_mem_counter[1042] = 4'b0000;
    GSharePlugin_logic_mem_counter[1043] = 4'b0000;
    GSharePlugin_logic_mem_counter[1044] = 4'b0000;
    GSharePlugin_logic_mem_counter[1045] = 4'b0000;
    GSharePlugin_logic_mem_counter[1046] = 4'b0000;
    GSharePlugin_logic_mem_counter[1047] = 4'b0000;
    GSharePlugin_logic_mem_counter[1048] = 4'b0000;
    GSharePlugin_logic_mem_counter[1049] = 4'b0000;
    GSharePlugin_logic_mem_counter[1050] = 4'b0000;
    GSharePlugin_logic_mem_counter[1051] = 4'b0000;
    GSharePlugin_logic_mem_counter[1052] = 4'b0000;
    GSharePlugin_logic_mem_counter[1053] = 4'b0000;
    GSharePlugin_logic_mem_counter[1054] = 4'b0000;
    GSharePlugin_logic_mem_counter[1055] = 4'b0000;
    GSharePlugin_logic_mem_counter[1056] = 4'b0000;
    GSharePlugin_logic_mem_counter[1057] = 4'b0000;
    GSharePlugin_logic_mem_counter[1058] = 4'b0000;
    GSharePlugin_logic_mem_counter[1059] = 4'b0000;
    GSharePlugin_logic_mem_counter[1060] = 4'b0000;
    GSharePlugin_logic_mem_counter[1061] = 4'b0000;
    GSharePlugin_logic_mem_counter[1062] = 4'b0000;
    GSharePlugin_logic_mem_counter[1063] = 4'b0000;
    GSharePlugin_logic_mem_counter[1064] = 4'b0000;
    GSharePlugin_logic_mem_counter[1065] = 4'b0000;
    GSharePlugin_logic_mem_counter[1066] = 4'b0000;
    GSharePlugin_logic_mem_counter[1067] = 4'b0000;
    GSharePlugin_logic_mem_counter[1068] = 4'b0000;
    GSharePlugin_logic_mem_counter[1069] = 4'b0000;
    GSharePlugin_logic_mem_counter[1070] = 4'b0000;
    GSharePlugin_logic_mem_counter[1071] = 4'b0000;
    GSharePlugin_logic_mem_counter[1072] = 4'b0000;
    GSharePlugin_logic_mem_counter[1073] = 4'b0000;
    GSharePlugin_logic_mem_counter[1074] = 4'b0000;
    GSharePlugin_logic_mem_counter[1075] = 4'b0000;
    GSharePlugin_logic_mem_counter[1076] = 4'b0000;
    GSharePlugin_logic_mem_counter[1077] = 4'b0000;
    GSharePlugin_logic_mem_counter[1078] = 4'b0000;
    GSharePlugin_logic_mem_counter[1079] = 4'b0000;
    GSharePlugin_logic_mem_counter[1080] = 4'b0000;
    GSharePlugin_logic_mem_counter[1081] = 4'b0000;
    GSharePlugin_logic_mem_counter[1082] = 4'b0000;
    GSharePlugin_logic_mem_counter[1083] = 4'b0000;
    GSharePlugin_logic_mem_counter[1084] = 4'b0000;
    GSharePlugin_logic_mem_counter[1085] = 4'b0000;
    GSharePlugin_logic_mem_counter[1086] = 4'b0000;
    GSharePlugin_logic_mem_counter[1087] = 4'b0000;
    GSharePlugin_logic_mem_counter[1088] = 4'b0000;
    GSharePlugin_logic_mem_counter[1089] = 4'b0000;
    GSharePlugin_logic_mem_counter[1090] = 4'b0000;
    GSharePlugin_logic_mem_counter[1091] = 4'b0000;
    GSharePlugin_logic_mem_counter[1092] = 4'b0000;
    GSharePlugin_logic_mem_counter[1093] = 4'b0000;
    GSharePlugin_logic_mem_counter[1094] = 4'b0000;
    GSharePlugin_logic_mem_counter[1095] = 4'b0000;
    GSharePlugin_logic_mem_counter[1096] = 4'b0000;
    GSharePlugin_logic_mem_counter[1097] = 4'b0000;
    GSharePlugin_logic_mem_counter[1098] = 4'b0000;
    GSharePlugin_logic_mem_counter[1099] = 4'b0000;
    GSharePlugin_logic_mem_counter[1100] = 4'b0000;
    GSharePlugin_logic_mem_counter[1101] = 4'b0000;
    GSharePlugin_logic_mem_counter[1102] = 4'b0000;
    GSharePlugin_logic_mem_counter[1103] = 4'b0000;
    GSharePlugin_logic_mem_counter[1104] = 4'b0000;
    GSharePlugin_logic_mem_counter[1105] = 4'b0000;
    GSharePlugin_logic_mem_counter[1106] = 4'b0000;
    GSharePlugin_logic_mem_counter[1107] = 4'b0000;
    GSharePlugin_logic_mem_counter[1108] = 4'b0000;
    GSharePlugin_logic_mem_counter[1109] = 4'b0000;
    GSharePlugin_logic_mem_counter[1110] = 4'b0000;
    GSharePlugin_logic_mem_counter[1111] = 4'b0000;
    GSharePlugin_logic_mem_counter[1112] = 4'b0000;
    GSharePlugin_logic_mem_counter[1113] = 4'b0000;
    GSharePlugin_logic_mem_counter[1114] = 4'b0000;
    GSharePlugin_logic_mem_counter[1115] = 4'b0000;
    GSharePlugin_logic_mem_counter[1116] = 4'b0000;
    GSharePlugin_logic_mem_counter[1117] = 4'b0000;
    GSharePlugin_logic_mem_counter[1118] = 4'b0000;
    GSharePlugin_logic_mem_counter[1119] = 4'b0000;
    GSharePlugin_logic_mem_counter[1120] = 4'b0000;
    GSharePlugin_logic_mem_counter[1121] = 4'b0000;
    GSharePlugin_logic_mem_counter[1122] = 4'b0000;
    GSharePlugin_logic_mem_counter[1123] = 4'b0000;
    GSharePlugin_logic_mem_counter[1124] = 4'b0000;
    GSharePlugin_logic_mem_counter[1125] = 4'b0000;
    GSharePlugin_logic_mem_counter[1126] = 4'b0000;
    GSharePlugin_logic_mem_counter[1127] = 4'b0000;
    GSharePlugin_logic_mem_counter[1128] = 4'b0000;
    GSharePlugin_logic_mem_counter[1129] = 4'b0000;
    GSharePlugin_logic_mem_counter[1130] = 4'b0000;
    GSharePlugin_logic_mem_counter[1131] = 4'b0000;
    GSharePlugin_logic_mem_counter[1132] = 4'b0000;
    GSharePlugin_logic_mem_counter[1133] = 4'b0000;
    GSharePlugin_logic_mem_counter[1134] = 4'b0000;
    GSharePlugin_logic_mem_counter[1135] = 4'b0000;
    GSharePlugin_logic_mem_counter[1136] = 4'b0000;
    GSharePlugin_logic_mem_counter[1137] = 4'b0000;
    GSharePlugin_logic_mem_counter[1138] = 4'b0000;
    GSharePlugin_logic_mem_counter[1139] = 4'b0000;
    GSharePlugin_logic_mem_counter[1140] = 4'b0000;
    GSharePlugin_logic_mem_counter[1141] = 4'b0000;
    GSharePlugin_logic_mem_counter[1142] = 4'b0000;
    GSharePlugin_logic_mem_counter[1143] = 4'b0000;
    GSharePlugin_logic_mem_counter[1144] = 4'b0000;
    GSharePlugin_logic_mem_counter[1145] = 4'b0000;
    GSharePlugin_logic_mem_counter[1146] = 4'b0000;
    GSharePlugin_logic_mem_counter[1147] = 4'b0000;
    GSharePlugin_logic_mem_counter[1148] = 4'b0000;
    GSharePlugin_logic_mem_counter[1149] = 4'b0000;
    GSharePlugin_logic_mem_counter[1150] = 4'b0000;
    GSharePlugin_logic_mem_counter[1151] = 4'b0000;
    GSharePlugin_logic_mem_counter[1152] = 4'b0000;
    GSharePlugin_logic_mem_counter[1153] = 4'b0000;
    GSharePlugin_logic_mem_counter[1154] = 4'b0000;
    GSharePlugin_logic_mem_counter[1155] = 4'b0000;
    GSharePlugin_logic_mem_counter[1156] = 4'b0000;
    GSharePlugin_logic_mem_counter[1157] = 4'b0000;
    GSharePlugin_logic_mem_counter[1158] = 4'b0000;
    GSharePlugin_logic_mem_counter[1159] = 4'b0000;
    GSharePlugin_logic_mem_counter[1160] = 4'b0000;
    GSharePlugin_logic_mem_counter[1161] = 4'b0000;
    GSharePlugin_logic_mem_counter[1162] = 4'b0000;
    GSharePlugin_logic_mem_counter[1163] = 4'b0000;
    GSharePlugin_logic_mem_counter[1164] = 4'b0000;
    GSharePlugin_logic_mem_counter[1165] = 4'b0000;
    GSharePlugin_logic_mem_counter[1166] = 4'b0000;
    GSharePlugin_logic_mem_counter[1167] = 4'b0000;
    GSharePlugin_logic_mem_counter[1168] = 4'b0000;
    GSharePlugin_logic_mem_counter[1169] = 4'b0000;
    GSharePlugin_logic_mem_counter[1170] = 4'b0000;
    GSharePlugin_logic_mem_counter[1171] = 4'b0000;
    GSharePlugin_logic_mem_counter[1172] = 4'b0000;
    GSharePlugin_logic_mem_counter[1173] = 4'b0000;
    GSharePlugin_logic_mem_counter[1174] = 4'b0000;
    GSharePlugin_logic_mem_counter[1175] = 4'b0000;
    GSharePlugin_logic_mem_counter[1176] = 4'b0000;
    GSharePlugin_logic_mem_counter[1177] = 4'b0000;
    GSharePlugin_logic_mem_counter[1178] = 4'b0000;
    GSharePlugin_logic_mem_counter[1179] = 4'b0000;
    GSharePlugin_logic_mem_counter[1180] = 4'b0000;
    GSharePlugin_logic_mem_counter[1181] = 4'b0000;
    GSharePlugin_logic_mem_counter[1182] = 4'b0000;
    GSharePlugin_logic_mem_counter[1183] = 4'b0000;
    GSharePlugin_logic_mem_counter[1184] = 4'b0000;
    GSharePlugin_logic_mem_counter[1185] = 4'b0000;
    GSharePlugin_logic_mem_counter[1186] = 4'b0000;
    GSharePlugin_logic_mem_counter[1187] = 4'b0000;
    GSharePlugin_logic_mem_counter[1188] = 4'b0000;
    GSharePlugin_logic_mem_counter[1189] = 4'b0000;
    GSharePlugin_logic_mem_counter[1190] = 4'b0000;
    GSharePlugin_logic_mem_counter[1191] = 4'b0000;
    GSharePlugin_logic_mem_counter[1192] = 4'b0000;
    GSharePlugin_logic_mem_counter[1193] = 4'b0000;
    GSharePlugin_logic_mem_counter[1194] = 4'b0000;
    GSharePlugin_logic_mem_counter[1195] = 4'b0000;
    GSharePlugin_logic_mem_counter[1196] = 4'b0000;
    GSharePlugin_logic_mem_counter[1197] = 4'b0000;
    GSharePlugin_logic_mem_counter[1198] = 4'b0000;
    GSharePlugin_logic_mem_counter[1199] = 4'b0000;
    GSharePlugin_logic_mem_counter[1200] = 4'b0000;
    GSharePlugin_logic_mem_counter[1201] = 4'b0000;
    GSharePlugin_logic_mem_counter[1202] = 4'b0000;
    GSharePlugin_logic_mem_counter[1203] = 4'b0000;
    GSharePlugin_logic_mem_counter[1204] = 4'b0000;
    GSharePlugin_logic_mem_counter[1205] = 4'b0000;
    GSharePlugin_logic_mem_counter[1206] = 4'b0000;
    GSharePlugin_logic_mem_counter[1207] = 4'b0000;
    GSharePlugin_logic_mem_counter[1208] = 4'b0000;
    GSharePlugin_logic_mem_counter[1209] = 4'b0000;
    GSharePlugin_logic_mem_counter[1210] = 4'b0000;
    GSharePlugin_logic_mem_counter[1211] = 4'b0000;
    GSharePlugin_logic_mem_counter[1212] = 4'b0000;
    GSharePlugin_logic_mem_counter[1213] = 4'b0000;
    GSharePlugin_logic_mem_counter[1214] = 4'b0000;
    GSharePlugin_logic_mem_counter[1215] = 4'b0000;
    GSharePlugin_logic_mem_counter[1216] = 4'b0000;
    GSharePlugin_logic_mem_counter[1217] = 4'b0000;
    GSharePlugin_logic_mem_counter[1218] = 4'b0000;
    GSharePlugin_logic_mem_counter[1219] = 4'b0000;
    GSharePlugin_logic_mem_counter[1220] = 4'b0000;
    GSharePlugin_logic_mem_counter[1221] = 4'b0000;
    GSharePlugin_logic_mem_counter[1222] = 4'b0000;
    GSharePlugin_logic_mem_counter[1223] = 4'b0000;
    GSharePlugin_logic_mem_counter[1224] = 4'b0000;
    GSharePlugin_logic_mem_counter[1225] = 4'b0000;
    GSharePlugin_logic_mem_counter[1226] = 4'b0000;
    GSharePlugin_logic_mem_counter[1227] = 4'b0000;
    GSharePlugin_logic_mem_counter[1228] = 4'b0000;
    GSharePlugin_logic_mem_counter[1229] = 4'b0000;
    GSharePlugin_logic_mem_counter[1230] = 4'b0000;
    GSharePlugin_logic_mem_counter[1231] = 4'b0000;
    GSharePlugin_logic_mem_counter[1232] = 4'b0000;
    GSharePlugin_logic_mem_counter[1233] = 4'b0000;
    GSharePlugin_logic_mem_counter[1234] = 4'b0000;
    GSharePlugin_logic_mem_counter[1235] = 4'b0000;
    GSharePlugin_logic_mem_counter[1236] = 4'b0000;
    GSharePlugin_logic_mem_counter[1237] = 4'b0000;
    GSharePlugin_logic_mem_counter[1238] = 4'b0000;
    GSharePlugin_logic_mem_counter[1239] = 4'b0000;
    GSharePlugin_logic_mem_counter[1240] = 4'b0000;
    GSharePlugin_logic_mem_counter[1241] = 4'b0000;
    GSharePlugin_logic_mem_counter[1242] = 4'b0000;
    GSharePlugin_logic_mem_counter[1243] = 4'b0000;
    GSharePlugin_logic_mem_counter[1244] = 4'b0000;
    GSharePlugin_logic_mem_counter[1245] = 4'b0000;
    GSharePlugin_logic_mem_counter[1246] = 4'b0000;
    GSharePlugin_logic_mem_counter[1247] = 4'b0000;
    GSharePlugin_logic_mem_counter[1248] = 4'b0000;
    GSharePlugin_logic_mem_counter[1249] = 4'b0000;
    GSharePlugin_logic_mem_counter[1250] = 4'b0000;
    GSharePlugin_logic_mem_counter[1251] = 4'b0000;
    GSharePlugin_logic_mem_counter[1252] = 4'b0000;
    GSharePlugin_logic_mem_counter[1253] = 4'b0000;
    GSharePlugin_logic_mem_counter[1254] = 4'b0000;
    GSharePlugin_logic_mem_counter[1255] = 4'b0000;
    GSharePlugin_logic_mem_counter[1256] = 4'b0000;
    GSharePlugin_logic_mem_counter[1257] = 4'b0000;
    GSharePlugin_logic_mem_counter[1258] = 4'b0000;
    GSharePlugin_logic_mem_counter[1259] = 4'b0000;
    GSharePlugin_logic_mem_counter[1260] = 4'b0000;
    GSharePlugin_logic_mem_counter[1261] = 4'b0000;
    GSharePlugin_logic_mem_counter[1262] = 4'b0000;
    GSharePlugin_logic_mem_counter[1263] = 4'b0000;
    GSharePlugin_logic_mem_counter[1264] = 4'b0000;
    GSharePlugin_logic_mem_counter[1265] = 4'b0000;
    GSharePlugin_logic_mem_counter[1266] = 4'b0000;
    GSharePlugin_logic_mem_counter[1267] = 4'b0000;
    GSharePlugin_logic_mem_counter[1268] = 4'b0000;
    GSharePlugin_logic_mem_counter[1269] = 4'b0000;
    GSharePlugin_logic_mem_counter[1270] = 4'b0000;
    GSharePlugin_logic_mem_counter[1271] = 4'b0000;
    GSharePlugin_logic_mem_counter[1272] = 4'b0000;
    GSharePlugin_logic_mem_counter[1273] = 4'b0000;
    GSharePlugin_logic_mem_counter[1274] = 4'b0000;
    GSharePlugin_logic_mem_counter[1275] = 4'b0000;
    GSharePlugin_logic_mem_counter[1276] = 4'b0000;
    GSharePlugin_logic_mem_counter[1277] = 4'b0000;
    GSharePlugin_logic_mem_counter[1278] = 4'b0000;
    GSharePlugin_logic_mem_counter[1279] = 4'b0000;
    GSharePlugin_logic_mem_counter[1280] = 4'b0000;
    GSharePlugin_logic_mem_counter[1281] = 4'b0000;
    GSharePlugin_logic_mem_counter[1282] = 4'b0000;
    GSharePlugin_logic_mem_counter[1283] = 4'b0000;
    GSharePlugin_logic_mem_counter[1284] = 4'b0000;
    GSharePlugin_logic_mem_counter[1285] = 4'b0000;
    GSharePlugin_logic_mem_counter[1286] = 4'b0000;
    GSharePlugin_logic_mem_counter[1287] = 4'b0000;
    GSharePlugin_logic_mem_counter[1288] = 4'b0000;
    GSharePlugin_logic_mem_counter[1289] = 4'b0000;
    GSharePlugin_logic_mem_counter[1290] = 4'b0000;
    GSharePlugin_logic_mem_counter[1291] = 4'b0000;
    GSharePlugin_logic_mem_counter[1292] = 4'b0000;
    GSharePlugin_logic_mem_counter[1293] = 4'b0000;
    GSharePlugin_logic_mem_counter[1294] = 4'b0000;
    GSharePlugin_logic_mem_counter[1295] = 4'b0000;
    GSharePlugin_logic_mem_counter[1296] = 4'b0000;
    GSharePlugin_logic_mem_counter[1297] = 4'b0000;
    GSharePlugin_logic_mem_counter[1298] = 4'b0000;
    GSharePlugin_logic_mem_counter[1299] = 4'b0000;
    GSharePlugin_logic_mem_counter[1300] = 4'b0000;
    GSharePlugin_logic_mem_counter[1301] = 4'b0000;
    GSharePlugin_logic_mem_counter[1302] = 4'b0000;
    GSharePlugin_logic_mem_counter[1303] = 4'b0000;
    GSharePlugin_logic_mem_counter[1304] = 4'b0000;
    GSharePlugin_logic_mem_counter[1305] = 4'b0000;
    GSharePlugin_logic_mem_counter[1306] = 4'b0000;
    GSharePlugin_logic_mem_counter[1307] = 4'b0000;
    GSharePlugin_logic_mem_counter[1308] = 4'b0000;
    GSharePlugin_logic_mem_counter[1309] = 4'b0000;
    GSharePlugin_logic_mem_counter[1310] = 4'b0000;
    GSharePlugin_logic_mem_counter[1311] = 4'b0000;
    GSharePlugin_logic_mem_counter[1312] = 4'b0000;
    GSharePlugin_logic_mem_counter[1313] = 4'b0000;
    GSharePlugin_logic_mem_counter[1314] = 4'b0000;
    GSharePlugin_logic_mem_counter[1315] = 4'b0000;
    GSharePlugin_logic_mem_counter[1316] = 4'b0000;
    GSharePlugin_logic_mem_counter[1317] = 4'b0000;
    GSharePlugin_logic_mem_counter[1318] = 4'b0000;
    GSharePlugin_logic_mem_counter[1319] = 4'b0000;
    GSharePlugin_logic_mem_counter[1320] = 4'b0000;
    GSharePlugin_logic_mem_counter[1321] = 4'b0000;
    GSharePlugin_logic_mem_counter[1322] = 4'b0000;
    GSharePlugin_logic_mem_counter[1323] = 4'b0000;
    GSharePlugin_logic_mem_counter[1324] = 4'b0000;
    GSharePlugin_logic_mem_counter[1325] = 4'b0000;
    GSharePlugin_logic_mem_counter[1326] = 4'b0000;
    GSharePlugin_logic_mem_counter[1327] = 4'b0000;
    GSharePlugin_logic_mem_counter[1328] = 4'b0000;
    GSharePlugin_logic_mem_counter[1329] = 4'b0000;
    GSharePlugin_logic_mem_counter[1330] = 4'b0000;
    GSharePlugin_logic_mem_counter[1331] = 4'b0000;
    GSharePlugin_logic_mem_counter[1332] = 4'b0000;
    GSharePlugin_logic_mem_counter[1333] = 4'b0000;
    GSharePlugin_logic_mem_counter[1334] = 4'b0000;
    GSharePlugin_logic_mem_counter[1335] = 4'b0000;
    GSharePlugin_logic_mem_counter[1336] = 4'b0000;
    GSharePlugin_logic_mem_counter[1337] = 4'b0000;
    GSharePlugin_logic_mem_counter[1338] = 4'b0000;
    GSharePlugin_logic_mem_counter[1339] = 4'b0000;
    GSharePlugin_logic_mem_counter[1340] = 4'b0000;
    GSharePlugin_logic_mem_counter[1341] = 4'b0000;
    GSharePlugin_logic_mem_counter[1342] = 4'b0000;
    GSharePlugin_logic_mem_counter[1343] = 4'b0000;
    GSharePlugin_logic_mem_counter[1344] = 4'b0000;
    GSharePlugin_logic_mem_counter[1345] = 4'b0000;
    GSharePlugin_logic_mem_counter[1346] = 4'b0000;
    GSharePlugin_logic_mem_counter[1347] = 4'b0000;
    GSharePlugin_logic_mem_counter[1348] = 4'b0000;
    GSharePlugin_logic_mem_counter[1349] = 4'b0000;
    GSharePlugin_logic_mem_counter[1350] = 4'b0000;
    GSharePlugin_logic_mem_counter[1351] = 4'b0000;
    GSharePlugin_logic_mem_counter[1352] = 4'b0000;
    GSharePlugin_logic_mem_counter[1353] = 4'b0000;
    GSharePlugin_logic_mem_counter[1354] = 4'b0000;
    GSharePlugin_logic_mem_counter[1355] = 4'b0000;
    GSharePlugin_logic_mem_counter[1356] = 4'b0000;
    GSharePlugin_logic_mem_counter[1357] = 4'b0000;
    GSharePlugin_logic_mem_counter[1358] = 4'b0000;
    GSharePlugin_logic_mem_counter[1359] = 4'b0000;
    GSharePlugin_logic_mem_counter[1360] = 4'b0000;
    GSharePlugin_logic_mem_counter[1361] = 4'b0000;
    GSharePlugin_logic_mem_counter[1362] = 4'b0000;
    GSharePlugin_logic_mem_counter[1363] = 4'b0000;
    GSharePlugin_logic_mem_counter[1364] = 4'b0000;
    GSharePlugin_logic_mem_counter[1365] = 4'b0000;
    GSharePlugin_logic_mem_counter[1366] = 4'b0000;
    GSharePlugin_logic_mem_counter[1367] = 4'b0000;
    GSharePlugin_logic_mem_counter[1368] = 4'b0000;
    GSharePlugin_logic_mem_counter[1369] = 4'b0000;
    GSharePlugin_logic_mem_counter[1370] = 4'b0000;
    GSharePlugin_logic_mem_counter[1371] = 4'b0000;
    GSharePlugin_logic_mem_counter[1372] = 4'b0000;
    GSharePlugin_logic_mem_counter[1373] = 4'b0000;
    GSharePlugin_logic_mem_counter[1374] = 4'b0000;
    GSharePlugin_logic_mem_counter[1375] = 4'b0000;
    GSharePlugin_logic_mem_counter[1376] = 4'b0000;
    GSharePlugin_logic_mem_counter[1377] = 4'b0000;
    GSharePlugin_logic_mem_counter[1378] = 4'b0000;
    GSharePlugin_logic_mem_counter[1379] = 4'b0000;
    GSharePlugin_logic_mem_counter[1380] = 4'b0000;
    GSharePlugin_logic_mem_counter[1381] = 4'b0000;
    GSharePlugin_logic_mem_counter[1382] = 4'b0000;
    GSharePlugin_logic_mem_counter[1383] = 4'b0000;
    GSharePlugin_logic_mem_counter[1384] = 4'b0000;
    GSharePlugin_logic_mem_counter[1385] = 4'b0000;
    GSharePlugin_logic_mem_counter[1386] = 4'b0000;
    GSharePlugin_logic_mem_counter[1387] = 4'b0000;
    GSharePlugin_logic_mem_counter[1388] = 4'b0000;
    GSharePlugin_logic_mem_counter[1389] = 4'b0000;
    GSharePlugin_logic_mem_counter[1390] = 4'b0000;
    GSharePlugin_logic_mem_counter[1391] = 4'b0000;
    GSharePlugin_logic_mem_counter[1392] = 4'b0000;
    GSharePlugin_logic_mem_counter[1393] = 4'b0000;
    GSharePlugin_logic_mem_counter[1394] = 4'b0000;
    GSharePlugin_logic_mem_counter[1395] = 4'b0000;
    GSharePlugin_logic_mem_counter[1396] = 4'b0000;
    GSharePlugin_logic_mem_counter[1397] = 4'b0000;
    GSharePlugin_logic_mem_counter[1398] = 4'b0000;
    GSharePlugin_logic_mem_counter[1399] = 4'b0000;
    GSharePlugin_logic_mem_counter[1400] = 4'b0000;
    GSharePlugin_logic_mem_counter[1401] = 4'b0000;
    GSharePlugin_logic_mem_counter[1402] = 4'b0000;
    GSharePlugin_logic_mem_counter[1403] = 4'b0000;
    GSharePlugin_logic_mem_counter[1404] = 4'b0000;
    GSharePlugin_logic_mem_counter[1405] = 4'b0000;
    GSharePlugin_logic_mem_counter[1406] = 4'b0000;
    GSharePlugin_logic_mem_counter[1407] = 4'b0000;
    GSharePlugin_logic_mem_counter[1408] = 4'b0000;
    GSharePlugin_logic_mem_counter[1409] = 4'b0000;
    GSharePlugin_logic_mem_counter[1410] = 4'b0000;
    GSharePlugin_logic_mem_counter[1411] = 4'b0000;
    GSharePlugin_logic_mem_counter[1412] = 4'b0000;
    GSharePlugin_logic_mem_counter[1413] = 4'b0000;
    GSharePlugin_logic_mem_counter[1414] = 4'b0000;
    GSharePlugin_logic_mem_counter[1415] = 4'b0000;
    GSharePlugin_logic_mem_counter[1416] = 4'b0000;
    GSharePlugin_logic_mem_counter[1417] = 4'b0000;
    GSharePlugin_logic_mem_counter[1418] = 4'b0000;
    GSharePlugin_logic_mem_counter[1419] = 4'b0000;
    GSharePlugin_logic_mem_counter[1420] = 4'b0000;
    GSharePlugin_logic_mem_counter[1421] = 4'b0000;
    GSharePlugin_logic_mem_counter[1422] = 4'b0000;
    GSharePlugin_logic_mem_counter[1423] = 4'b0000;
    GSharePlugin_logic_mem_counter[1424] = 4'b0000;
    GSharePlugin_logic_mem_counter[1425] = 4'b0000;
    GSharePlugin_logic_mem_counter[1426] = 4'b0000;
    GSharePlugin_logic_mem_counter[1427] = 4'b0000;
    GSharePlugin_logic_mem_counter[1428] = 4'b0000;
    GSharePlugin_logic_mem_counter[1429] = 4'b0000;
    GSharePlugin_logic_mem_counter[1430] = 4'b0000;
    GSharePlugin_logic_mem_counter[1431] = 4'b0000;
    GSharePlugin_logic_mem_counter[1432] = 4'b0000;
    GSharePlugin_logic_mem_counter[1433] = 4'b0000;
    GSharePlugin_logic_mem_counter[1434] = 4'b0000;
    GSharePlugin_logic_mem_counter[1435] = 4'b0000;
    GSharePlugin_logic_mem_counter[1436] = 4'b0000;
    GSharePlugin_logic_mem_counter[1437] = 4'b0000;
    GSharePlugin_logic_mem_counter[1438] = 4'b0000;
    GSharePlugin_logic_mem_counter[1439] = 4'b0000;
    GSharePlugin_logic_mem_counter[1440] = 4'b0000;
    GSharePlugin_logic_mem_counter[1441] = 4'b0000;
    GSharePlugin_logic_mem_counter[1442] = 4'b0000;
    GSharePlugin_logic_mem_counter[1443] = 4'b0000;
    GSharePlugin_logic_mem_counter[1444] = 4'b0000;
    GSharePlugin_logic_mem_counter[1445] = 4'b0000;
    GSharePlugin_logic_mem_counter[1446] = 4'b0000;
    GSharePlugin_logic_mem_counter[1447] = 4'b0000;
    GSharePlugin_logic_mem_counter[1448] = 4'b0000;
    GSharePlugin_logic_mem_counter[1449] = 4'b0000;
    GSharePlugin_logic_mem_counter[1450] = 4'b0000;
    GSharePlugin_logic_mem_counter[1451] = 4'b0000;
    GSharePlugin_logic_mem_counter[1452] = 4'b0000;
    GSharePlugin_logic_mem_counter[1453] = 4'b0000;
    GSharePlugin_logic_mem_counter[1454] = 4'b0000;
    GSharePlugin_logic_mem_counter[1455] = 4'b0000;
    GSharePlugin_logic_mem_counter[1456] = 4'b0000;
    GSharePlugin_logic_mem_counter[1457] = 4'b0000;
    GSharePlugin_logic_mem_counter[1458] = 4'b0000;
    GSharePlugin_logic_mem_counter[1459] = 4'b0000;
    GSharePlugin_logic_mem_counter[1460] = 4'b0000;
    GSharePlugin_logic_mem_counter[1461] = 4'b0000;
    GSharePlugin_logic_mem_counter[1462] = 4'b0000;
    GSharePlugin_logic_mem_counter[1463] = 4'b0000;
    GSharePlugin_logic_mem_counter[1464] = 4'b0000;
    GSharePlugin_logic_mem_counter[1465] = 4'b0000;
    GSharePlugin_logic_mem_counter[1466] = 4'b0000;
    GSharePlugin_logic_mem_counter[1467] = 4'b0000;
    GSharePlugin_logic_mem_counter[1468] = 4'b0000;
    GSharePlugin_logic_mem_counter[1469] = 4'b0000;
    GSharePlugin_logic_mem_counter[1470] = 4'b0000;
    GSharePlugin_logic_mem_counter[1471] = 4'b0000;
    GSharePlugin_logic_mem_counter[1472] = 4'b0000;
    GSharePlugin_logic_mem_counter[1473] = 4'b0000;
    GSharePlugin_logic_mem_counter[1474] = 4'b0000;
    GSharePlugin_logic_mem_counter[1475] = 4'b0000;
    GSharePlugin_logic_mem_counter[1476] = 4'b0000;
    GSharePlugin_logic_mem_counter[1477] = 4'b0000;
    GSharePlugin_logic_mem_counter[1478] = 4'b0000;
    GSharePlugin_logic_mem_counter[1479] = 4'b0000;
    GSharePlugin_logic_mem_counter[1480] = 4'b0000;
    GSharePlugin_logic_mem_counter[1481] = 4'b0000;
    GSharePlugin_logic_mem_counter[1482] = 4'b0000;
    GSharePlugin_logic_mem_counter[1483] = 4'b0000;
    GSharePlugin_logic_mem_counter[1484] = 4'b0000;
    GSharePlugin_logic_mem_counter[1485] = 4'b0000;
    GSharePlugin_logic_mem_counter[1486] = 4'b0000;
    GSharePlugin_logic_mem_counter[1487] = 4'b0000;
    GSharePlugin_logic_mem_counter[1488] = 4'b0000;
    GSharePlugin_logic_mem_counter[1489] = 4'b0000;
    GSharePlugin_logic_mem_counter[1490] = 4'b0000;
    GSharePlugin_logic_mem_counter[1491] = 4'b0000;
    GSharePlugin_logic_mem_counter[1492] = 4'b0000;
    GSharePlugin_logic_mem_counter[1493] = 4'b0000;
    GSharePlugin_logic_mem_counter[1494] = 4'b0000;
    GSharePlugin_logic_mem_counter[1495] = 4'b0000;
    GSharePlugin_logic_mem_counter[1496] = 4'b0000;
    GSharePlugin_logic_mem_counter[1497] = 4'b0000;
    GSharePlugin_logic_mem_counter[1498] = 4'b0000;
    GSharePlugin_logic_mem_counter[1499] = 4'b0000;
    GSharePlugin_logic_mem_counter[1500] = 4'b0000;
    GSharePlugin_logic_mem_counter[1501] = 4'b0000;
    GSharePlugin_logic_mem_counter[1502] = 4'b0000;
    GSharePlugin_logic_mem_counter[1503] = 4'b0000;
    GSharePlugin_logic_mem_counter[1504] = 4'b0000;
    GSharePlugin_logic_mem_counter[1505] = 4'b0000;
    GSharePlugin_logic_mem_counter[1506] = 4'b0000;
    GSharePlugin_logic_mem_counter[1507] = 4'b0000;
    GSharePlugin_logic_mem_counter[1508] = 4'b0000;
    GSharePlugin_logic_mem_counter[1509] = 4'b0000;
    GSharePlugin_logic_mem_counter[1510] = 4'b0000;
    GSharePlugin_logic_mem_counter[1511] = 4'b0000;
    GSharePlugin_logic_mem_counter[1512] = 4'b0000;
    GSharePlugin_logic_mem_counter[1513] = 4'b0000;
    GSharePlugin_logic_mem_counter[1514] = 4'b0000;
    GSharePlugin_logic_mem_counter[1515] = 4'b0000;
    GSharePlugin_logic_mem_counter[1516] = 4'b0000;
    GSharePlugin_logic_mem_counter[1517] = 4'b0000;
    GSharePlugin_logic_mem_counter[1518] = 4'b0000;
    GSharePlugin_logic_mem_counter[1519] = 4'b0000;
    GSharePlugin_logic_mem_counter[1520] = 4'b0000;
    GSharePlugin_logic_mem_counter[1521] = 4'b0000;
    GSharePlugin_logic_mem_counter[1522] = 4'b0000;
    GSharePlugin_logic_mem_counter[1523] = 4'b0000;
    GSharePlugin_logic_mem_counter[1524] = 4'b0000;
    GSharePlugin_logic_mem_counter[1525] = 4'b0000;
    GSharePlugin_logic_mem_counter[1526] = 4'b0000;
    GSharePlugin_logic_mem_counter[1527] = 4'b0000;
    GSharePlugin_logic_mem_counter[1528] = 4'b0000;
    GSharePlugin_logic_mem_counter[1529] = 4'b0000;
    GSharePlugin_logic_mem_counter[1530] = 4'b0000;
    GSharePlugin_logic_mem_counter[1531] = 4'b0000;
    GSharePlugin_logic_mem_counter[1532] = 4'b0000;
    GSharePlugin_logic_mem_counter[1533] = 4'b0000;
    GSharePlugin_logic_mem_counter[1534] = 4'b0000;
    GSharePlugin_logic_mem_counter[1535] = 4'b0000;
    GSharePlugin_logic_mem_counter[1536] = 4'b0000;
    GSharePlugin_logic_mem_counter[1537] = 4'b0000;
    GSharePlugin_logic_mem_counter[1538] = 4'b0000;
    GSharePlugin_logic_mem_counter[1539] = 4'b0000;
    GSharePlugin_logic_mem_counter[1540] = 4'b0000;
    GSharePlugin_logic_mem_counter[1541] = 4'b0000;
    GSharePlugin_logic_mem_counter[1542] = 4'b0000;
    GSharePlugin_logic_mem_counter[1543] = 4'b0000;
    GSharePlugin_logic_mem_counter[1544] = 4'b0000;
    GSharePlugin_logic_mem_counter[1545] = 4'b0000;
    GSharePlugin_logic_mem_counter[1546] = 4'b0000;
    GSharePlugin_logic_mem_counter[1547] = 4'b0000;
    GSharePlugin_logic_mem_counter[1548] = 4'b0000;
    GSharePlugin_logic_mem_counter[1549] = 4'b0000;
    GSharePlugin_logic_mem_counter[1550] = 4'b0000;
    GSharePlugin_logic_mem_counter[1551] = 4'b0000;
    GSharePlugin_logic_mem_counter[1552] = 4'b0000;
    GSharePlugin_logic_mem_counter[1553] = 4'b0000;
    GSharePlugin_logic_mem_counter[1554] = 4'b0000;
    GSharePlugin_logic_mem_counter[1555] = 4'b0000;
    GSharePlugin_logic_mem_counter[1556] = 4'b0000;
    GSharePlugin_logic_mem_counter[1557] = 4'b0000;
    GSharePlugin_logic_mem_counter[1558] = 4'b0000;
    GSharePlugin_logic_mem_counter[1559] = 4'b0000;
    GSharePlugin_logic_mem_counter[1560] = 4'b0000;
    GSharePlugin_logic_mem_counter[1561] = 4'b0000;
    GSharePlugin_logic_mem_counter[1562] = 4'b0000;
    GSharePlugin_logic_mem_counter[1563] = 4'b0000;
    GSharePlugin_logic_mem_counter[1564] = 4'b0000;
    GSharePlugin_logic_mem_counter[1565] = 4'b0000;
    GSharePlugin_logic_mem_counter[1566] = 4'b0000;
    GSharePlugin_logic_mem_counter[1567] = 4'b0000;
    GSharePlugin_logic_mem_counter[1568] = 4'b0000;
    GSharePlugin_logic_mem_counter[1569] = 4'b0000;
    GSharePlugin_logic_mem_counter[1570] = 4'b0000;
    GSharePlugin_logic_mem_counter[1571] = 4'b0000;
    GSharePlugin_logic_mem_counter[1572] = 4'b0000;
    GSharePlugin_logic_mem_counter[1573] = 4'b0000;
    GSharePlugin_logic_mem_counter[1574] = 4'b0000;
    GSharePlugin_logic_mem_counter[1575] = 4'b0000;
    GSharePlugin_logic_mem_counter[1576] = 4'b0000;
    GSharePlugin_logic_mem_counter[1577] = 4'b0000;
    GSharePlugin_logic_mem_counter[1578] = 4'b0000;
    GSharePlugin_logic_mem_counter[1579] = 4'b0000;
    GSharePlugin_logic_mem_counter[1580] = 4'b0000;
    GSharePlugin_logic_mem_counter[1581] = 4'b0000;
    GSharePlugin_logic_mem_counter[1582] = 4'b0000;
    GSharePlugin_logic_mem_counter[1583] = 4'b0000;
    GSharePlugin_logic_mem_counter[1584] = 4'b0000;
    GSharePlugin_logic_mem_counter[1585] = 4'b0000;
    GSharePlugin_logic_mem_counter[1586] = 4'b0000;
    GSharePlugin_logic_mem_counter[1587] = 4'b0000;
    GSharePlugin_logic_mem_counter[1588] = 4'b0000;
    GSharePlugin_logic_mem_counter[1589] = 4'b0000;
    GSharePlugin_logic_mem_counter[1590] = 4'b0000;
    GSharePlugin_logic_mem_counter[1591] = 4'b0000;
    GSharePlugin_logic_mem_counter[1592] = 4'b0000;
    GSharePlugin_logic_mem_counter[1593] = 4'b0000;
    GSharePlugin_logic_mem_counter[1594] = 4'b0000;
    GSharePlugin_logic_mem_counter[1595] = 4'b0000;
    GSharePlugin_logic_mem_counter[1596] = 4'b0000;
    GSharePlugin_logic_mem_counter[1597] = 4'b0000;
    GSharePlugin_logic_mem_counter[1598] = 4'b0000;
    GSharePlugin_logic_mem_counter[1599] = 4'b0000;
    GSharePlugin_logic_mem_counter[1600] = 4'b0000;
    GSharePlugin_logic_mem_counter[1601] = 4'b0000;
    GSharePlugin_logic_mem_counter[1602] = 4'b0000;
    GSharePlugin_logic_mem_counter[1603] = 4'b0000;
    GSharePlugin_logic_mem_counter[1604] = 4'b0000;
    GSharePlugin_logic_mem_counter[1605] = 4'b0000;
    GSharePlugin_logic_mem_counter[1606] = 4'b0000;
    GSharePlugin_logic_mem_counter[1607] = 4'b0000;
    GSharePlugin_logic_mem_counter[1608] = 4'b0000;
    GSharePlugin_logic_mem_counter[1609] = 4'b0000;
    GSharePlugin_logic_mem_counter[1610] = 4'b0000;
    GSharePlugin_logic_mem_counter[1611] = 4'b0000;
    GSharePlugin_logic_mem_counter[1612] = 4'b0000;
    GSharePlugin_logic_mem_counter[1613] = 4'b0000;
    GSharePlugin_logic_mem_counter[1614] = 4'b0000;
    GSharePlugin_logic_mem_counter[1615] = 4'b0000;
    GSharePlugin_logic_mem_counter[1616] = 4'b0000;
    GSharePlugin_logic_mem_counter[1617] = 4'b0000;
    GSharePlugin_logic_mem_counter[1618] = 4'b0000;
    GSharePlugin_logic_mem_counter[1619] = 4'b0000;
    GSharePlugin_logic_mem_counter[1620] = 4'b0000;
    GSharePlugin_logic_mem_counter[1621] = 4'b0000;
    GSharePlugin_logic_mem_counter[1622] = 4'b0000;
    GSharePlugin_logic_mem_counter[1623] = 4'b0000;
    GSharePlugin_logic_mem_counter[1624] = 4'b0000;
    GSharePlugin_logic_mem_counter[1625] = 4'b0000;
    GSharePlugin_logic_mem_counter[1626] = 4'b0000;
    GSharePlugin_logic_mem_counter[1627] = 4'b0000;
    GSharePlugin_logic_mem_counter[1628] = 4'b0000;
    GSharePlugin_logic_mem_counter[1629] = 4'b0000;
    GSharePlugin_logic_mem_counter[1630] = 4'b0000;
    GSharePlugin_logic_mem_counter[1631] = 4'b0000;
    GSharePlugin_logic_mem_counter[1632] = 4'b0000;
    GSharePlugin_logic_mem_counter[1633] = 4'b0000;
    GSharePlugin_logic_mem_counter[1634] = 4'b0000;
    GSharePlugin_logic_mem_counter[1635] = 4'b0000;
    GSharePlugin_logic_mem_counter[1636] = 4'b0000;
    GSharePlugin_logic_mem_counter[1637] = 4'b0000;
    GSharePlugin_logic_mem_counter[1638] = 4'b0000;
    GSharePlugin_logic_mem_counter[1639] = 4'b0000;
    GSharePlugin_logic_mem_counter[1640] = 4'b0000;
    GSharePlugin_logic_mem_counter[1641] = 4'b0000;
    GSharePlugin_logic_mem_counter[1642] = 4'b0000;
    GSharePlugin_logic_mem_counter[1643] = 4'b0000;
    GSharePlugin_logic_mem_counter[1644] = 4'b0000;
    GSharePlugin_logic_mem_counter[1645] = 4'b0000;
    GSharePlugin_logic_mem_counter[1646] = 4'b0000;
    GSharePlugin_logic_mem_counter[1647] = 4'b0000;
    GSharePlugin_logic_mem_counter[1648] = 4'b0000;
    GSharePlugin_logic_mem_counter[1649] = 4'b0000;
    GSharePlugin_logic_mem_counter[1650] = 4'b0000;
    GSharePlugin_logic_mem_counter[1651] = 4'b0000;
    GSharePlugin_logic_mem_counter[1652] = 4'b0000;
    GSharePlugin_logic_mem_counter[1653] = 4'b0000;
    GSharePlugin_logic_mem_counter[1654] = 4'b0000;
    GSharePlugin_logic_mem_counter[1655] = 4'b0000;
    GSharePlugin_logic_mem_counter[1656] = 4'b0000;
    GSharePlugin_logic_mem_counter[1657] = 4'b0000;
    GSharePlugin_logic_mem_counter[1658] = 4'b0000;
    GSharePlugin_logic_mem_counter[1659] = 4'b0000;
    GSharePlugin_logic_mem_counter[1660] = 4'b0000;
    GSharePlugin_logic_mem_counter[1661] = 4'b0000;
    GSharePlugin_logic_mem_counter[1662] = 4'b0000;
    GSharePlugin_logic_mem_counter[1663] = 4'b0000;
    GSharePlugin_logic_mem_counter[1664] = 4'b0000;
    GSharePlugin_logic_mem_counter[1665] = 4'b0000;
    GSharePlugin_logic_mem_counter[1666] = 4'b0000;
    GSharePlugin_logic_mem_counter[1667] = 4'b0000;
    GSharePlugin_logic_mem_counter[1668] = 4'b0000;
    GSharePlugin_logic_mem_counter[1669] = 4'b0000;
    GSharePlugin_logic_mem_counter[1670] = 4'b0000;
    GSharePlugin_logic_mem_counter[1671] = 4'b0000;
    GSharePlugin_logic_mem_counter[1672] = 4'b0000;
    GSharePlugin_logic_mem_counter[1673] = 4'b0000;
    GSharePlugin_logic_mem_counter[1674] = 4'b0000;
    GSharePlugin_logic_mem_counter[1675] = 4'b0000;
    GSharePlugin_logic_mem_counter[1676] = 4'b0000;
    GSharePlugin_logic_mem_counter[1677] = 4'b0000;
    GSharePlugin_logic_mem_counter[1678] = 4'b0000;
    GSharePlugin_logic_mem_counter[1679] = 4'b0000;
    GSharePlugin_logic_mem_counter[1680] = 4'b0000;
    GSharePlugin_logic_mem_counter[1681] = 4'b0000;
    GSharePlugin_logic_mem_counter[1682] = 4'b0000;
    GSharePlugin_logic_mem_counter[1683] = 4'b0000;
    GSharePlugin_logic_mem_counter[1684] = 4'b0000;
    GSharePlugin_logic_mem_counter[1685] = 4'b0000;
    GSharePlugin_logic_mem_counter[1686] = 4'b0000;
    GSharePlugin_logic_mem_counter[1687] = 4'b0000;
    GSharePlugin_logic_mem_counter[1688] = 4'b0000;
    GSharePlugin_logic_mem_counter[1689] = 4'b0000;
    GSharePlugin_logic_mem_counter[1690] = 4'b0000;
    GSharePlugin_logic_mem_counter[1691] = 4'b0000;
    GSharePlugin_logic_mem_counter[1692] = 4'b0000;
    GSharePlugin_logic_mem_counter[1693] = 4'b0000;
    GSharePlugin_logic_mem_counter[1694] = 4'b0000;
    GSharePlugin_logic_mem_counter[1695] = 4'b0000;
    GSharePlugin_logic_mem_counter[1696] = 4'b0000;
    GSharePlugin_logic_mem_counter[1697] = 4'b0000;
    GSharePlugin_logic_mem_counter[1698] = 4'b0000;
    GSharePlugin_logic_mem_counter[1699] = 4'b0000;
    GSharePlugin_logic_mem_counter[1700] = 4'b0000;
    GSharePlugin_logic_mem_counter[1701] = 4'b0000;
    GSharePlugin_logic_mem_counter[1702] = 4'b0000;
    GSharePlugin_logic_mem_counter[1703] = 4'b0000;
    GSharePlugin_logic_mem_counter[1704] = 4'b0000;
    GSharePlugin_logic_mem_counter[1705] = 4'b0000;
    GSharePlugin_logic_mem_counter[1706] = 4'b0000;
    GSharePlugin_logic_mem_counter[1707] = 4'b0000;
    GSharePlugin_logic_mem_counter[1708] = 4'b0000;
    GSharePlugin_logic_mem_counter[1709] = 4'b0000;
    GSharePlugin_logic_mem_counter[1710] = 4'b0000;
    GSharePlugin_logic_mem_counter[1711] = 4'b0000;
    GSharePlugin_logic_mem_counter[1712] = 4'b0000;
    GSharePlugin_logic_mem_counter[1713] = 4'b0000;
    GSharePlugin_logic_mem_counter[1714] = 4'b0000;
    GSharePlugin_logic_mem_counter[1715] = 4'b0000;
    GSharePlugin_logic_mem_counter[1716] = 4'b0000;
    GSharePlugin_logic_mem_counter[1717] = 4'b0000;
    GSharePlugin_logic_mem_counter[1718] = 4'b0000;
    GSharePlugin_logic_mem_counter[1719] = 4'b0000;
    GSharePlugin_logic_mem_counter[1720] = 4'b0000;
    GSharePlugin_logic_mem_counter[1721] = 4'b0000;
    GSharePlugin_logic_mem_counter[1722] = 4'b0000;
    GSharePlugin_logic_mem_counter[1723] = 4'b0000;
    GSharePlugin_logic_mem_counter[1724] = 4'b0000;
    GSharePlugin_logic_mem_counter[1725] = 4'b0000;
    GSharePlugin_logic_mem_counter[1726] = 4'b0000;
    GSharePlugin_logic_mem_counter[1727] = 4'b0000;
    GSharePlugin_logic_mem_counter[1728] = 4'b0000;
    GSharePlugin_logic_mem_counter[1729] = 4'b0000;
    GSharePlugin_logic_mem_counter[1730] = 4'b0000;
    GSharePlugin_logic_mem_counter[1731] = 4'b0000;
    GSharePlugin_logic_mem_counter[1732] = 4'b0000;
    GSharePlugin_logic_mem_counter[1733] = 4'b0000;
    GSharePlugin_logic_mem_counter[1734] = 4'b0000;
    GSharePlugin_logic_mem_counter[1735] = 4'b0000;
    GSharePlugin_logic_mem_counter[1736] = 4'b0000;
    GSharePlugin_logic_mem_counter[1737] = 4'b0000;
    GSharePlugin_logic_mem_counter[1738] = 4'b0000;
    GSharePlugin_logic_mem_counter[1739] = 4'b0000;
    GSharePlugin_logic_mem_counter[1740] = 4'b0000;
    GSharePlugin_logic_mem_counter[1741] = 4'b0000;
    GSharePlugin_logic_mem_counter[1742] = 4'b0000;
    GSharePlugin_logic_mem_counter[1743] = 4'b0000;
    GSharePlugin_logic_mem_counter[1744] = 4'b0000;
    GSharePlugin_logic_mem_counter[1745] = 4'b0000;
    GSharePlugin_logic_mem_counter[1746] = 4'b0000;
    GSharePlugin_logic_mem_counter[1747] = 4'b0000;
    GSharePlugin_logic_mem_counter[1748] = 4'b0000;
    GSharePlugin_logic_mem_counter[1749] = 4'b0000;
    GSharePlugin_logic_mem_counter[1750] = 4'b0000;
    GSharePlugin_logic_mem_counter[1751] = 4'b0000;
    GSharePlugin_logic_mem_counter[1752] = 4'b0000;
    GSharePlugin_logic_mem_counter[1753] = 4'b0000;
    GSharePlugin_logic_mem_counter[1754] = 4'b0000;
    GSharePlugin_logic_mem_counter[1755] = 4'b0000;
    GSharePlugin_logic_mem_counter[1756] = 4'b0000;
    GSharePlugin_logic_mem_counter[1757] = 4'b0000;
    GSharePlugin_logic_mem_counter[1758] = 4'b0000;
    GSharePlugin_logic_mem_counter[1759] = 4'b0000;
    GSharePlugin_logic_mem_counter[1760] = 4'b0000;
    GSharePlugin_logic_mem_counter[1761] = 4'b0000;
    GSharePlugin_logic_mem_counter[1762] = 4'b0000;
    GSharePlugin_logic_mem_counter[1763] = 4'b0000;
    GSharePlugin_logic_mem_counter[1764] = 4'b0000;
    GSharePlugin_logic_mem_counter[1765] = 4'b0000;
    GSharePlugin_logic_mem_counter[1766] = 4'b0000;
    GSharePlugin_logic_mem_counter[1767] = 4'b0000;
    GSharePlugin_logic_mem_counter[1768] = 4'b0000;
    GSharePlugin_logic_mem_counter[1769] = 4'b0000;
    GSharePlugin_logic_mem_counter[1770] = 4'b0000;
    GSharePlugin_logic_mem_counter[1771] = 4'b0000;
    GSharePlugin_logic_mem_counter[1772] = 4'b0000;
    GSharePlugin_logic_mem_counter[1773] = 4'b0000;
    GSharePlugin_logic_mem_counter[1774] = 4'b0000;
    GSharePlugin_logic_mem_counter[1775] = 4'b0000;
    GSharePlugin_logic_mem_counter[1776] = 4'b0000;
    GSharePlugin_logic_mem_counter[1777] = 4'b0000;
    GSharePlugin_logic_mem_counter[1778] = 4'b0000;
    GSharePlugin_logic_mem_counter[1779] = 4'b0000;
    GSharePlugin_logic_mem_counter[1780] = 4'b0000;
    GSharePlugin_logic_mem_counter[1781] = 4'b0000;
    GSharePlugin_logic_mem_counter[1782] = 4'b0000;
    GSharePlugin_logic_mem_counter[1783] = 4'b0000;
    GSharePlugin_logic_mem_counter[1784] = 4'b0000;
    GSharePlugin_logic_mem_counter[1785] = 4'b0000;
    GSharePlugin_logic_mem_counter[1786] = 4'b0000;
    GSharePlugin_logic_mem_counter[1787] = 4'b0000;
    GSharePlugin_logic_mem_counter[1788] = 4'b0000;
    GSharePlugin_logic_mem_counter[1789] = 4'b0000;
    GSharePlugin_logic_mem_counter[1790] = 4'b0000;
    GSharePlugin_logic_mem_counter[1791] = 4'b0000;
    GSharePlugin_logic_mem_counter[1792] = 4'b0000;
    GSharePlugin_logic_mem_counter[1793] = 4'b0000;
    GSharePlugin_logic_mem_counter[1794] = 4'b0000;
    GSharePlugin_logic_mem_counter[1795] = 4'b0000;
    GSharePlugin_logic_mem_counter[1796] = 4'b0000;
    GSharePlugin_logic_mem_counter[1797] = 4'b0000;
    GSharePlugin_logic_mem_counter[1798] = 4'b0000;
    GSharePlugin_logic_mem_counter[1799] = 4'b0000;
    GSharePlugin_logic_mem_counter[1800] = 4'b0000;
    GSharePlugin_logic_mem_counter[1801] = 4'b0000;
    GSharePlugin_logic_mem_counter[1802] = 4'b0000;
    GSharePlugin_logic_mem_counter[1803] = 4'b0000;
    GSharePlugin_logic_mem_counter[1804] = 4'b0000;
    GSharePlugin_logic_mem_counter[1805] = 4'b0000;
    GSharePlugin_logic_mem_counter[1806] = 4'b0000;
    GSharePlugin_logic_mem_counter[1807] = 4'b0000;
    GSharePlugin_logic_mem_counter[1808] = 4'b0000;
    GSharePlugin_logic_mem_counter[1809] = 4'b0000;
    GSharePlugin_logic_mem_counter[1810] = 4'b0000;
    GSharePlugin_logic_mem_counter[1811] = 4'b0000;
    GSharePlugin_logic_mem_counter[1812] = 4'b0000;
    GSharePlugin_logic_mem_counter[1813] = 4'b0000;
    GSharePlugin_logic_mem_counter[1814] = 4'b0000;
    GSharePlugin_logic_mem_counter[1815] = 4'b0000;
    GSharePlugin_logic_mem_counter[1816] = 4'b0000;
    GSharePlugin_logic_mem_counter[1817] = 4'b0000;
    GSharePlugin_logic_mem_counter[1818] = 4'b0000;
    GSharePlugin_logic_mem_counter[1819] = 4'b0000;
    GSharePlugin_logic_mem_counter[1820] = 4'b0000;
    GSharePlugin_logic_mem_counter[1821] = 4'b0000;
    GSharePlugin_logic_mem_counter[1822] = 4'b0000;
    GSharePlugin_logic_mem_counter[1823] = 4'b0000;
    GSharePlugin_logic_mem_counter[1824] = 4'b0000;
    GSharePlugin_logic_mem_counter[1825] = 4'b0000;
    GSharePlugin_logic_mem_counter[1826] = 4'b0000;
    GSharePlugin_logic_mem_counter[1827] = 4'b0000;
    GSharePlugin_logic_mem_counter[1828] = 4'b0000;
    GSharePlugin_logic_mem_counter[1829] = 4'b0000;
    GSharePlugin_logic_mem_counter[1830] = 4'b0000;
    GSharePlugin_logic_mem_counter[1831] = 4'b0000;
    GSharePlugin_logic_mem_counter[1832] = 4'b0000;
    GSharePlugin_logic_mem_counter[1833] = 4'b0000;
    GSharePlugin_logic_mem_counter[1834] = 4'b0000;
    GSharePlugin_logic_mem_counter[1835] = 4'b0000;
    GSharePlugin_logic_mem_counter[1836] = 4'b0000;
    GSharePlugin_logic_mem_counter[1837] = 4'b0000;
    GSharePlugin_logic_mem_counter[1838] = 4'b0000;
    GSharePlugin_logic_mem_counter[1839] = 4'b0000;
    GSharePlugin_logic_mem_counter[1840] = 4'b0000;
    GSharePlugin_logic_mem_counter[1841] = 4'b0000;
    GSharePlugin_logic_mem_counter[1842] = 4'b0000;
    GSharePlugin_logic_mem_counter[1843] = 4'b0000;
    GSharePlugin_logic_mem_counter[1844] = 4'b0000;
    GSharePlugin_logic_mem_counter[1845] = 4'b0000;
    GSharePlugin_logic_mem_counter[1846] = 4'b0000;
    GSharePlugin_logic_mem_counter[1847] = 4'b0000;
    GSharePlugin_logic_mem_counter[1848] = 4'b0000;
    GSharePlugin_logic_mem_counter[1849] = 4'b0000;
    GSharePlugin_logic_mem_counter[1850] = 4'b0000;
    GSharePlugin_logic_mem_counter[1851] = 4'b0000;
    GSharePlugin_logic_mem_counter[1852] = 4'b0000;
    GSharePlugin_logic_mem_counter[1853] = 4'b0000;
    GSharePlugin_logic_mem_counter[1854] = 4'b0000;
    GSharePlugin_logic_mem_counter[1855] = 4'b0000;
    GSharePlugin_logic_mem_counter[1856] = 4'b0000;
    GSharePlugin_logic_mem_counter[1857] = 4'b0000;
    GSharePlugin_logic_mem_counter[1858] = 4'b0000;
    GSharePlugin_logic_mem_counter[1859] = 4'b0000;
    GSharePlugin_logic_mem_counter[1860] = 4'b0000;
    GSharePlugin_logic_mem_counter[1861] = 4'b0000;
    GSharePlugin_logic_mem_counter[1862] = 4'b0000;
    GSharePlugin_logic_mem_counter[1863] = 4'b0000;
    GSharePlugin_logic_mem_counter[1864] = 4'b0000;
    GSharePlugin_logic_mem_counter[1865] = 4'b0000;
    GSharePlugin_logic_mem_counter[1866] = 4'b0000;
    GSharePlugin_logic_mem_counter[1867] = 4'b0000;
    GSharePlugin_logic_mem_counter[1868] = 4'b0000;
    GSharePlugin_logic_mem_counter[1869] = 4'b0000;
    GSharePlugin_logic_mem_counter[1870] = 4'b0000;
    GSharePlugin_logic_mem_counter[1871] = 4'b0000;
    GSharePlugin_logic_mem_counter[1872] = 4'b0000;
    GSharePlugin_logic_mem_counter[1873] = 4'b0000;
    GSharePlugin_logic_mem_counter[1874] = 4'b0000;
    GSharePlugin_logic_mem_counter[1875] = 4'b0000;
    GSharePlugin_logic_mem_counter[1876] = 4'b0000;
    GSharePlugin_logic_mem_counter[1877] = 4'b0000;
    GSharePlugin_logic_mem_counter[1878] = 4'b0000;
    GSharePlugin_logic_mem_counter[1879] = 4'b0000;
    GSharePlugin_logic_mem_counter[1880] = 4'b0000;
    GSharePlugin_logic_mem_counter[1881] = 4'b0000;
    GSharePlugin_logic_mem_counter[1882] = 4'b0000;
    GSharePlugin_logic_mem_counter[1883] = 4'b0000;
    GSharePlugin_logic_mem_counter[1884] = 4'b0000;
    GSharePlugin_logic_mem_counter[1885] = 4'b0000;
    GSharePlugin_logic_mem_counter[1886] = 4'b0000;
    GSharePlugin_logic_mem_counter[1887] = 4'b0000;
    GSharePlugin_logic_mem_counter[1888] = 4'b0000;
    GSharePlugin_logic_mem_counter[1889] = 4'b0000;
    GSharePlugin_logic_mem_counter[1890] = 4'b0000;
    GSharePlugin_logic_mem_counter[1891] = 4'b0000;
    GSharePlugin_logic_mem_counter[1892] = 4'b0000;
    GSharePlugin_logic_mem_counter[1893] = 4'b0000;
    GSharePlugin_logic_mem_counter[1894] = 4'b0000;
    GSharePlugin_logic_mem_counter[1895] = 4'b0000;
    GSharePlugin_logic_mem_counter[1896] = 4'b0000;
    GSharePlugin_logic_mem_counter[1897] = 4'b0000;
    GSharePlugin_logic_mem_counter[1898] = 4'b0000;
    GSharePlugin_logic_mem_counter[1899] = 4'b0000;
    GSharePlugin_logic_mem_counter[1900] = 4'b0000;
    GSharePlugin_logic_mem_counter[1901] = 4'b0000;
    GSharePlugin_logic_mem_counter[1902] = 4'b0000;
    GSharePlugin_logic_mem_counter[1903] = 4'b0000;
    GSharePlugin_logic_mem_counter[1904] = 4'b0000;
    GSharePlugin_logic_mem_counter[1905] = 4'b0000;
    GSharePlugin_logic_mem_counter[1906] = 4'b0000;
    GSharePlugin_logic_mem_counter[1907] = 4'b0000;
    GSharePlugin_logic_mem_counter[1908] = 4'b0000;
    GSharePlugin_logic_mem_counter[1909] = 4'b0000;
    GSharePlugin_logic_mem_counter[1910] = 4'b0000;
    GSharePlugin_logic_mem_counter[1911] = 4'b0000;
    GSharePlugin_logic_mem_counter[1912] = 4'b0000;
    GSharePlugin_logic_mem_counter[1913] = 4'b0000;
    GSharePlugin_logic_mem_counter[1914] = 4'b0000;
    GSharePlugin_logic_mem_counter[1915] = 4'b0000;
    GSharePlugin_logic_mem_counter[1916] = 4'b0000;
    GSharePlugin_logic_mem_counter[1917] = 4'b0000;
    GSharePlugin_logic_mem_counter[1918] = 4'b0000;
    GSharePlugin_logic_mem_counter[1919] = 4'b0000;
    GSharePlugin_logic_mem_counter[1920] = 4'b0000;
    GSharePlugin_logic_mem_counter[1921] = 4'b0000;
    GSharePlugin_logic_mem_counter[1922] = 4'b0000;
    GSharePlugin_logic_mem_counter[1923] = 4'b0000;
    GSharePlugin_logic_mem_counter[1924] = 4'b0000;
    GSharePlugin_logic_mem_counter[1925] = 4'b0000;
    GSharePlugin_logic_mem_counter[1926] = 4'b0000;
    GSharePlugin_logic_mem_counter[1927] = 4'b0000;
    GSharePlugin_logic_mem_counter[1928] = 4'b0000;
    GSharePlugin_logic_mem_counter[1929] = 4'b0000;
    GSharePlugin_logic_mem_counter[1930] = 4'b0000;
    GSharePlugin_logic_mem_counter[1931] = 4'b0000;
    GSharePlugin_logic_mem_counter[1932] = 4'b0000;
    GSharePlugin_logic_mem_counter[1933] = 4'b0000;
    GSharePlugin_logic_mem_counter[1934] = 4'b0000;
    GSharePlugin_logic_mem_counter[1935] = 4'b0000;
    GSharePlugin_logic_mem_counter[1936] = 4'b0000;
    GSharePlugin_logic_mem_counter[1937] = 4'b0000;
    GSharePlugin_logic_mem_counter[1938] = 4'b0000;
    GSharePlugin_logic_mem_counter[1939] = 4'b0000;
    GSharePlugin_logic_mem_counter[1940] = 4'b0000;
    GSharePlugin_logic_mem_counter[1941] = 4'b0000;
    GSharePlugin_logic_mem_counter[1942] = 4'b0000;
    GSharePlugin_logic_mem_counter[1943] = 4'b0000;
    GSharePlugin_logic_mem_counter[1944] = 4'b0000;
    GSharePlugin_logic_mem_counter[1945] = 4'b0000;
    GSharePlugin_logic_mem_counter[1946] = 4'b0000;
    GSharePlugin_logic_mem_counter[1947] = 4'b0000;
    GSharePlugin_logic_mem_counter[1948] = 4'b0000;
    GSharePlugin_logic_mem_counter[1949] = 4'b0000;
    GSharePlugin_logic_mem_counter[1950] = 4'b0000;
    GSharePlugin_logic_mem_counter[1951] = 4'b0000;
    GSharePlugin_logic_mem_counter[1952] = 4'b0000;
    GSharePlugin_logic_mem_counter[1953] = 4'b0000;
    GSharePlugin_logic_mem_counter[1954] = 4'b0000;
    GSharePlugin_logic_mem_counter[1955] = 4'b0000;
    GSharePlugin_logic_mem_counter[1956] = 4'b0000;
    GSharePlugin_logic_mem_counter[1957] = 4'b0000;
    GSharePlugin_logic_mem_counter[1958] = 4'b0000;
    GSharePlugin_logic_mem_counter[1959] = 4'b0000;
    GSharePlugin_logic_mem_counter[1960] = 4'b0000;
    GSharePlugin_logic_mem_counter[1961] = 4'b0000;
    GSharePlugin_logic_mem_counter[1962] = 4'b0000;
    GSharePlugin_logic_mem_counter[1963] = 4'b0000;
    GSharePlugin_logic_mem_counter[1964] = 4'b0000;
    GSharePlugin_logic_mem_counter[1965] = 4'b0000;
    GSharePlugin_logic_mem_counter[1966] = 4'b0000;
    GSharePlugin_logic_mem_counter[1967] = 4'b0000;
    GSharePlugin_logic_mem_counter[1968] = 4'b0000;
    GSharePlugin_logic_mem_counter[1969] = 4'b0000;
    GSharePlugin_logic_mem_counter[1970] = 4'b0000;
    GSharePlugin_logic_mem_counter[1971] = 4'b0000;
    GSharePlugin_logic_mem_counter[1972] = 4'b0000;
    GSharePlugin_logic_mem_counter[1973] = 4'b0000;
    GSharePlugin_logic_mem_counter[1974] = 4'b0000;
    GSharePlugin_logic_mem_counter[1975] = 4'b0000;
    GSharePlugin_logic_mem_counter[1976] = 4'b0000;
    GSharePlugin_logic_mem_counter[1977] = 4'b0000;
    GSharePlugin_logic_mem_counter[1978] = 4'b0000;
    GSharePlugin_logic_mem_counter[1979] = 4'b0000;
    GSharePlugin_logic_mem_counter[1980] = 4'b0000;
    GSharePlugin_logic_mem_counter[1981] = 4'b0000;
    GSharePlugin_logic_mem_counter[1982] = 4'b0000;
    GSharePlugin_logic_mem_counter[1983] = 4'b0000;
    GSharePlugin_logic_mem_counter[1984] = 4'b0000;
    GSharePlugin_logic_mem_counter[1985] = 4'b0000;
    GSharePlugin_logic_mem_counter[1986] = 4'b0000;
    GSharePlugin_logic_mem_counter[1987] = 4'b0000;
    GSharePlugin_logic_mem_counter[1988] = 4'b0000;
    GSharePlugin_logic_mem_counter[1989] = 4'b0000;
    GSharePlugin_logic_mem_counter[1990] = 4'b0000;
    GSharePlugin_logic_mem_counter[1991] = 4'b0000;
    GSharePlugin_logic_mem_counter[1992] = 4'b0000;
    GSharePlugin_logic_mem_counter[1993] = 4'b0000;
    GSharePlugin_logic_mem_counter[1994] = 4'b0000;
    GSharePlugin_logic_mem_counter[1995] = 4'b0000;
    GSharePlugin_logic_mem_counter[1996] = 4'b0000;
    GSharePlugin_logic_mem_counter[1997] = 4'b0000;
    GSharePlugin_logic_mem_counter[1998] = 4'b0000;
    GSharePlugin_logic_mem_counter[1999] = 4'b0000;
    GSharePlugin_logic_mem_counter[2000] = 4'b0000;
    GSharePlugin_logic_mem_counter[2001] = 4'b0000;
    GSharePlugin_logic_mem_counter[2002] = 4'b0000;
    GSharePlugin_logic_mem_counter[2003] = 4'b0000;
    GSharePlugin_logic_mem_counter[2004] = 4'b0000;
    GSharePlugin_logic_mem_counter[2005] = 4'b0000;
    GSharePlugin_logic_mem_counter[2006] = 4'b0000;
    GSharePlugin_logic_mem_counter[2007] = 4'b0000;
    GSharePlugin_logic_mem_counter[2008] = 4'b0000;
    GSharePlugin_logic_mem_counter[2009] = 4'b0000;
    GSharePlugin_logic_mem_counter[2010] = 4'b0000;
    GSharePlugin_logic_mem_counter[2011] = 4'b0000;
    GSharePlugin_logic_mem_counter[2012] = 4'b0000;
    GSharePlugin_logic_mem_counter[2013] = 4'b0000;
    GSharePlugin_logic_mem_counter[2014] = 4'b0000;
    GSharePlugin_logic_mem_counter[2015] = 4'b0000;
    GSharePlugin_logic_mem_counter[2016] = 4'b0000;
    GSharePlugin_logic_mem_counter[2017] = 4'b0000;
    GSharePlugin_logic_mem_counter[2018] = 4'b0000;
    GSharePlugin_logic_mem_counter[2019] = 4'b0000;
    GSharePlugin_logic_mem_counter[2020] = 4'b0000;
    GSharePlugin_logic_mem_counter[2021] = 4'b0000;
    GSharePlugin_logic_mem_counter[2022] = 4'b0000;
    GSharePlugin_logic_mem_counter[2023] = 4'b0000;
    GSharePlugin_logic_mem_counter[2024] = 4'b0000;
    GSharePlugin_logic_mem_counter[2025] = 4'b0000;
    GSharePlugin_logic_mem_counter[2026] = 4'b0000;
    GSharePlugin_logic_mem_counter[2027] = 4'b0000;
    GSharePlugin_logic_mem_counter[2028] = 4'b0000;
    GSharePlugin_logic_mem_counter[2029] = 4'b0000;
    GSharePlugin_logic_mem_counter[2030] = 4'b0000;
    GSharePlugin_logic_mem_counter[2031] = 4'b0000;
    GSharePlugin_logic_mem_counter[2032] = 4'b0000;
    GSharePlugin_logic_mem_counter[2033] = 4'b0000;
    GSharePlugin_logic_mem_counter[2034] = 4'b0000;
    GSharePlugin_logic_mem_counter[2035] = 4'b0000;
    GSharePlugin_logic_mem_counter[2036] = 4'b0000;
    GSharePlugin_logic_mem_counter[2037] = 4'b0000;
    GSharePlugin_logic_mem_counter[2038] = 4'b0000;
    GSharePlugin_logic_mem_counter[2039] = 4'b0000;
    GSharePlugin_logic_mem_counter[2040] = 4'b0000;
    GSharePlugin_logic_mem_counter[2041] = 4'b0000;
    GSharePlugin_logic_mem_counter[2042] = 4'b0000;
    GSharePlugin_logic_mem_counter[2043] = 4'b0000;
    GSharePlugin_logic_mem_counter[2044] = 4'b0000;
    GSharePlugin_logic_mem_counter[2045] = 4'b0000;
    GSharePlugin_logic_mem_counter[2046] = 4'b0000;
    GSharePlugin_logic_mem_counter[2047] = 4'b0000;
    GSharePlugin_logic_mem_counter[2048] = 4'b0000;
    GSharePlugin_logic_mem_counter[2049] = 4'b0000;
    GSharePlugin_logic_mem_counter[2050] = 4'b0000;
    GSharePlugin_logic_mem_counter[2051] = 4'b0000;
    GSharePlugin_logic_mem_counter[2052] = 4'b0000;
    GSharePlugin_logic_mem_counter[2053] = 4'b0000;
    GSharePlugin_logic_mem_counter[2054] = 4'b0000;
    GSharePlugin_logic_mem_counter[2055] = 4'b0000;
    GSharePlugin_logic_mem_counter[2056] = 4'b0000;
    GSharePlugin_logic_mem_counter[2057] = 4'b0000;
    GSharePlugin_logic_mem_counter[2058] = 4'b0000;
    GSharePlugin_logic_mem_counter[2059] = 4'b0000;
    GSharePlugin_logic_mem_counter[2060] = 4'b0000;
    GSharePlugin_logic_mem_counter[2061] = 4'b0000;
    GSharePlugin_logic_mem_counter[2062] = 4'b0000;
    GSharePlugin_logic_mem_counter[2063] = 4'b0000;
    GSharePlugin_logic_mem_counter[2064] = 4'b0000;
    GSharePlugin_logic_mem_counter[2065] = 4'b0000;
    GSharePlugin_logic_mem_counter[2066] = 4'b0000;
    GSharePlugin_logic_mem_counter[2067] = 4'b0000;
    GSharePlugin_logic_mem_counter[2068] = 4'b0000;
    GSharePlugin_logic_mem_counter[2069] = 4'b0000;
    GSharePlugin_logic_mem_counter[2070] = 4'b0000;
    GSharePlugin_logic_mem_counter[2071] = 4'b0000;
    GSharePlugin_logic_mem_counter[2072] = 4'b0000;
    GSharePlugin_logic_mem_counter[2073] = 4'b0000;
    GSharePlugin_logic_mem_counter[2074] = 4'b0000;
    GSharePlugin_logic_mem_counter[2075] = 4'b0000;
    GSharePlugin_logic_mem_counter[2076] = 4'b0000;
    GSharePlugin_logic_mem_counter[2077] = 4'b0000;
    GSharePlugin_logic_mem_counter[2078] = 4'b0000;
    GSharePlugin_logic_mem_counter[2079] = 4'b0000;
    GSharePlugin_logic_mem_counter[2080] = 4'b0000;
    GSharePlugin_logic_mem_counter[2081] = 4'b0000;
    GSharePlugin_logic_mem_counter[2082] = 4'b0000;
    GSharePlugin_logic_mem_counter[2083] = 4'b0000;
    GSharePlugin_logic_mem_counter[2084] = 4'b0000;
    GSharePlugin_logic_mem_counter[2085] = 4'b0000;
    GSharePlugin_logic_mem_counter[2086] = 4'b0000;
    GSharePlugin_logic_mem_counter[2087] = 4'b0000;
    GSharePlugin_logic_mem_counter[2088] = 4'b0000;
    GSharePlugin_logic_mem_counter[2089] = 4'b0000;
    GSharePlugin_logic_mem_counter[2090] = 4'b0000;
    GSharePlugin_logic_mem_counter[2091] = 4'b0000;
    GSharePlugin_logic_mem_counter[2092] = 4'b0000;
    GSharePlugin_logic_mem_counter[2093] = 4'b0000;
    GSharePlugin_logic_mem_counter[2094] = 4'b0000;
    GSharePlugin_logic_mem_counter[2095] = 4'b0000;
    GSharePlugin_logic_mem_counter[2096] = 4'b0000;
    GSharePlugin_logic_mem_counter[2097] = 4'b0000;
    GSharePlugin_logic_mem_counter[2098] = 4'b0000;
    GSharePlugin_logic_mem_counter[2099] = 4'b0000;
    GSharePlugin_logic_mem_counter[2100] = 4'b0000;
    GSharePlugin_logic_mem_counter[2101] = 4'b0000;
    GSharePlugin_logic_mem_counter[2102] = 4'b0000;
    GSharePlugin_logic_mem_counter[2103] = 4'b0000;
    GSharePlugin_logic_mem_counter[2104] = 4'b0000;
    GSharePlugin_logic_mem_counter[2105] = 4'b0000;
    GSharePlugin_logic_mem_counter[2106] = 4'b0000;
    GSharePlugin_logic_mem_counter[2107] = 4'b0000;
    GSharePlugin_logic_mem_counter[2108] = 4'b0000;
    GSharePlugin_logic_mem_counter[2109] = 4'b0000;
    GSharePlugin_logic_mem_counter[2110] = 4'b0000;
    GSharePlugin_logic_mem_counter[2111] = 4'b0000;
    GSharePlugin_logic_mem_counter[2112] = 4'b0000;
    GSharePlugin_logic_mem_counter[2113] = 4'b0000;
    GSharePlugin_logic_mem_counter[2114] = 4'b0000;
    GSharePlugin_logic_mem_counter[2115] = 4'b0000;
    GSharePlugin_logic_mem_counter[2116] = 4'b0000;
    GSharePlugin_logic_mem_counter[2117] = 4'b0000;
    GSharePlugin_logic_mem_counter[2118] = 4'b0000;
    GSharePlugin_logic_mem_counter[2119] = 4'b0000;
    GSharePlugin_logic_mem_counter[2120] = 4'b0000;
    GSharePlugin_logic_mem_counter[2121] = 4'b0000;
    GSharePlugin_logic_mem_counter[2122] = 4'b0000;
    GSharePlugin_logic_mem_counter[2123] = 4'b0000;
    GSharePlugin_logic_mem_counter[2124] = 4'b0000;
    GSharePlugin_logic_mem_counter[2125] = 4'b0000;
    GSharePlugin_logic_mem_counter[2126] = 4'b0000;
    GSharePlugin_logic_mem_counter[2127] = 4'b0000;
    GSharePlugin_logic_mem_counter[2128] = 4'b0000;
    GSharePlugin_logic_mem_counter[2129] = 4'b0000;
    GSharePlugin_logic_mem_counter[2130] = 4'b0000;
    GSharePlugin_logic_mem_counter[2131] = 4'b0000;
    GSharePlugin_logic_mem_counter[2132] = 4'b0000;
    GSharePlugin_logic_mem_counter[2133] = 4'b0000;
    GSharePlugin_logic_mem_counter[2134] = 4'b0000;
    GSharePlugin_logic_mem_counter[2135] = 4'b0000;
    GSharePlugin_logic_mem_counter[2136] = 4'b0000;
    GSharePlugin_logic_mem_counter[2137] = 4'b0000;
    GSharePlugin_logic_mem_counter[2138] = 4'b0000;
    GSharePlugin_logic_mem_counter[2139] = 4'b0000;
    GSharePlugin_logic_mem_counter[2140] = 4'b0000;
    GSharePlugin_logic_mem_counter[2141] = 4'b0000;
    GSharePlugin_logic_mem_counter[2142] = 4'b0000;
    GSharePlugin_logic_mem_counter[2143] = 4'b0000;
    GSharePlugin_logic_mem_counter[2144] = 4'b0000;
    GSharePlugin_logic_mem_counter[2145] = 4'b0000;
    GSharePlugin_logic_mem_counter[2146] = 4'b0000;
    GSharePlugin_logic_mem_counter[2147] = 4'b0000;
    GSharePlugin_logic_mem_counter[2148] = 4'b0000;
    GSharePlugin_logic_mem_counter[2149] = 4'b0000;
    GSharePlugin_logic_mem_counter[2150] = 4'b0000;
    GSharePlugin_logic_mem_counter[2151] = 4'b0000;
    GSharePlugin_logic_mem_counter[2152] = 4'b0000;
    GSharePlugin_logic_mem_counter[2153] = 4'b0000;
    GSharePlugin_logic_mem_counter[2154] = 4'b0000;
    GSharePlugin_logic_mem_counter[2155] = 4'b0000;
    GSharePlugin_logic_mem_counter[2156] = 4'b0000;
    GSharePlugin_logic_mem_counter[2157] = 4'b0000;
    GSharePlugin_logic_mem_counter[2158] = 4'b0000;
    GSharePlugin_logic_mem_counter[2159] = 4'b0000;
    GSharePlugin_logic_mem_counter[2160] = 4'b0000;
    GSharePlugin_logic_mem_counter[2161] = 4'b0000;
    GSharePlugin_logic_mem_counter[2162] = 4'b0000;
    GSharePlugin_logic_mem_counter[2163] = 4'b0000;
    GSharePlugin_logic_mem_counter[2164] = 4'b0000;
    GSharePlugin_logic_mem_counter[2165] = 4'b0000;
    GSharePlugin_logic_mem_counter[2166] = 4'b0000;
    GSharePlugin_logic_mem_counter[2167] = 4'b0000;
    GSharePlugin_logic_mem_counter[2168] = 4'b0000;
    GSharePlugin_logic_mem_counter[2169] = 4'b0000;
    GSharePlugin_logic_mem_counter[2170] = 4'b0000;
    GSharePlugin_logic_mem_counter[2171] = 4'b0000;
    GSharePlugin_logic_mem_counter[2172] = 4'b0000;
    GSharePlugin_logic_mem_counter[2173] = 4'b0000;
    GSharePlugin_logic_mem_counter[2174] = 4'b0000;
    GSharePlugin_logic_mem_counter[2175] = 4'b0000;
    GSharePlugin_logic_mem_counter[2176] = 4'b0000;
    GSharePlugin_logic_mem_counter[2177] = 4'b0000;
    GSharePlugin_logic_mem_counter[2178] = 4'b0000;
    GSharePlugin_logic_mem_counter[2179] = 4'b0000;
    GSharePlugin_logic_mem_counter[2180] = 4'b0000;
    GSharePlugin_logic_mem_counter[2181] = 4'b0000;
    GSharePlugin_logic_mem_counter[2182] = 4'b0000;
    GSharePlugin_logic_mem_counter[2183] = 4'b0000;
    GSharePlugin_logic_mem_counter[2184] = 4'b0000;
    GSharePlugin_logic_mem_counter[2185] = 4'b0000;
    GSharePlugin_logic_mem_counter[2186] = 4'b0000;
    GSharePlugin_logic_mem_counter[2187] = 4'b0000;
    GSharePlugin_logic_mem_counter[2188] = 4'b0000;
    GSharePlugin_logic_mem_counter[2189] = 4'b0000;
    GSharePlugin_logic_mem_counter[2190] = 4'b0000;
    GSharePlugin_logic_mem_counter[2191] = 4'b0000;
    GSharePlugin_logic_mem_counter[2192] = 4'b0000;
    GSharePlugin_logic_mem_counter[2193] = 4'b0000;
    GSharePlugin_logic_mem_counter[2194] = 4'b0000;
    GSharePlugin_logic_mem_counter[2195] = 4'b0000;
    GSharePlugin_logic_mem_counter[2196] = 4'b0000;
    GSharePlugin_logic_mem_counter[2197] = 4'b0000;
    GSharePlugin_logic_mem_counter[2198] = 4'b0000;
    GSharePlugin_logic_mem_counter[2199] = 4'b0000;
    GSharePlugin_logic_mem_counter[2200] = 4'b0000;
    GSharePlugin_logic_mem_counter[2201] = 4'b0000;
    GSharePlugin_logic_mem_counter[2202] = 4'b0000;
    GSharePlugin_logic_mem_counter[2203] = 4'b0000;
    GSharePlugin_logic_mem_counter[2204] = 4'b0000;
    GSharePlugin_logic_mem_counter[2205] = 4'b0000;
    GSharePlugin_logic_mem_counter[2206] = 4'b0000;
    GSharePlugin_logic_mem_counter[2207] = 4'b0000;
    GSharePlugin_logic_mem_counter[2208] = 4'b0000;
    GSharePlugin_logic_mem_counter[2209] = 4'b0000;
    GSharePlugin_logic_mem_counter[2210] = 4'b0000;
    GSharePlugin_logic_mem_counter[2211] = 4'b0000;
    GSharePlugin_logic_mem_counter[2212] = 4'b0000;
    GSharePlugin_logic_mem_counter[2213] = 4'b0000;
    GSharePlugin_logic_mem_counter[2214] = 4'b0000;
    GSharePlugin_logic_mem_counter[2215] = 4'b0000;
    GSharePlugin_logic_mem_counter[2216] = 4'b0000;
    GSharePlugin_logic_mem_counter[2217] = 4'b0000;
    GSharePlugin_logic_mem_counter[2218] = 4'b0000;
    GSharePlugin_logic_mem_counter[2219] = 4'b0000;
    GSharePlugin_logic_mem_counter[2220] = 4'b0000;
    GSharePlugin_logic_mem_counter[2221] = 4'b0000;
    GSharePlugin_logic_mem_counter[2222] = 4'b0000;
    GSharePlugin_logic_mem_counter[2223] = 4'b0000;
    GSharePlugin_logic_mem_counter[2224] = 4'b0000;
    GSharePlugin_logic_mem_counter[2225] = 4'b0000;
    GSharePlugin_logic_mem_counter[2226] = 4'b0000;
    GSharePlugin_logic_mem_counter[2227] = 4'b0000;
    GSharePlugin_logic_mem_counter[2228] = 4'b0000;
    GSharePlugin_logic_mem_counter[2229] = 4'b0000;
    GSharePlugin_logic_mem_counter[2230] = 4'b0000;
    GSharePlugin_logic_mem_counter[2231] = 4'b0000;
    GSharePlugin_logic_mem_counter[2232] = 4'b0000;
    GSharePlugin_logic_mem_counter[2233] = 4'b0000;
    GSharePlugin_logic_mem_counter[2234] = 4'b0000;
    GSharePlugin_logic_mem_counter[2235] = 4'b0000;
    GSharePlugin_logic_mem_counter[2236] = 4'b0000;
    GSharePlugin_logic_mem_counter[2237] = 4'b0000;
    GSharePlugin_logic_mem_counter[2238] = 4'b0000;
    GSharePlugin_logic_mem_counter[2239] = 4'b0000;
    GSharePlugin_logic_mem_counter[2240] = 4'b0000;
    GSharePlugin_logic_mem_counter[2241] = 4'b0000;
    GSharePlugin_logic_mem_counter[2242] = 4'b0000;
    GSharePlugin_logic_mem_counter[2243] = 4'b0000;
    GSharePlugin_logic_mem_counter[2244] = 4'b0000;
    GSharePlugin_logic_mem_counter[2245] = 4'b0000;
    GSharePlugin_logic_mem_counter[2246] = 4'b0000;
    GSharePlugin_logic_mem_counter[2247] = 4'b0000;
    GSharePlugin_logic_mem_counter[2248] = 4'b0000;
    GSharePlugin_logic_mem_counter[2249] = 4'b0000;
    GSharePlugin_logic_mem_counter[2250] = 4'b0000;
    GSharePlugin_logic_mem_counter[2251] = 4'b0000;
    GSharePlugin_logic_mem_counter[2252] = 4'b0000;
    GSharePlugin_logic_mem_counter[2253] = 4'b0000;
    GSharePlugin_logic_mem_counter[2254] = 4'b0000;
    GSharePlugin_logic_mem_counter[2255] = 4'b0000;
    GSharePlugin_logic_mem_counter[2256] = 4'b0000;
    GSharePlugin_logic_mem_counter[2257] = 4'b0000;
    GSharePlugin_logic_mem_counter[2258] = 4'b0000;
    GSharePlugin_logic_mem_counter[2259] = 4'b0000;
    GSharePlugin_logic_mem_counter[2260] = 4'b0000;
    GSharePlugin_logic_mem_counter[2261] = 4'b0000;
    GSharePlugin_logic_mem_counter[2262] = 4'b0000;
    GSharePlugin_logic_mem_counter[2263] = 4'b0000;
    GSharePlugin_logic_mem_counter[2264] = 4'b0000;
    GSharePlugin_logic_mem_counter[2265] = 4'b0000;
    GSharePlugin_logic_mem_counter[2266] = 4'b0000;
    GSharePlugin_logic_mem_counter[2267] = 4'b0000;
    GSharePlugin_logic_mem_counter[2268] = 4'b0000;
    GSharePlugin_logic_mem_counter[2269] = 4'b0000;
    GSharePlugin_logic_mem_counter[2270] = 4'b0000;
    GSharePlugin_logic_mem_counter[2271] = 4'b0000;
    GSharePlugin_logic_mem_counter[2272] = 4'b0000;
    GSharePlugin_logic_mem_counter[2273] = 4'b0000;
    GSharePlugin_logic_mem_counter[2274] = 4'b0000;
    GSharePlugin_logic_mem_counter[2275] = 4'b0000;
    GSharePlugin_logic_mem_counter[2276] = 4'b0000;
    GSharePlugin_logic_mem_counter[2277] = 4'b0000;
    GSharePlugin_logic_mem_counter[2278] = 4'b0000;
    GSharePlugin_logic_mem_counter[2279] = 4'b0000;
    GSharePlugin_logic_mem_counter[2280] = 4'b0000;
    GSharePlugin_logic_mem_counter[2281] = 4'b0000;
    GSharePlugin_logic_mem_counter[2282] = 4'b0000;
    GSharePlugin_logic_mem_counter[2283] = 4'b0000;
    GSharePlugin_logic_mem_counter[2284] = 4'b0000;
    GSharePlugin_logic_mem_counter[2285] = 4'b0000;
    GSharePlugin_logic_mem_counter[2286] = 4'b0000;
    GSharePlugin_logic_mem_counter[2287] = 4'b0000;
    GSharePlugin_logic_mem_counter[2288] = 4'b0000;
    GSharePlugin_logic_mem_counter[2289] = 4'b0000;
    GSharePlugin_logic_mem_counter[2290] = 4'b0000;
    GSharePlugin_logic_mem_counter[2291] = 4'b0000;
    GSharePlugin_logic_mem_counter[2292] = 4'b0000;
    GSharePlugin_logic_mem_counter[2293] = 4'b0000;
    GSharePlugin_logic_mem_counter[2294] = 4'b0000;
    GSharePlugin_logic_mem_counter[2295] = 4'b0000;
    GSharePlugin_logic_mem_counter[2296] = 4'b0000;
    GSharePlugin_logic_mem_counter[2297] = 4'b0000;
    GSharePlugin_logic_mem_counter[2298] = 4'b0000;
    GSharePlugin_logic_mem_counter[2299] = 4'b0000;
    GSharePlugin_logic_mem_counter[2300] = 4'b0000;
    GSharePlugin_logic_mem_counter[2301] = 4'b0000;
    GSharePlugin_logic_mem_counter[2302] = 4'b0000;
    GSharePlugin_logic_mem_counter[2303] = 4'b0000;
    GSharePlugin_logic_mem_counter[2304] = 4'b0000;
    GSharePlugin_logic_mem_counter[2305] = 4'b0000;
    GSharePlugin_logic_mem_counter[2306] = 4'b0000;
    GSharePlugin_logic_mem_counter[2307] = 4'b0000;
    GSharePlugin_logic_mem_counter[2308] = 4'b0000;
    GSharePlugin_logic_mem_counter[2309] = 4'b0000;
    GSharePlugin_logic_mem_counter[2310] = 4'b0000;
    GSharePlugin_logic_mem_counter[2311] = 4'b0000;
    GSharePlugin_logic_mem_counter[2312] = 4'b0000;
    GSharePlugin_logic_mem_counter[2313] = 4'b0000;
    GSharePlugin_logic_mem_counter[2314] = 4'b0000;
    GSharePlugin_logic_mem_counter[2315] = 4'b0000;
    GSharePlugin_logic_mem_counter[2316] = 4'b0000;
    GSharePlugin_logic_mem_counter[2317] = 4'b0000;
    GSharePlugin_logic_mem_counter[2318] = 4'b0000;
    GSharePlugin_logic_mem_counter[2319] = 4'b0000;
    GSharePlugin_logic_mem_counter[2320] = 4'b0000;
    GSharePlugin_logic_mem_counter[2321] = 4'b0000;
    GSharePlugin_logic_mem_counter[2322] = 4'b0000;
    GSharePlugin_logic_mem_counter[2323] = 4'b0000;
    GSharePlugin_logic_mem_counter[2324] = 4'b0000;
    GSharePlugin_logic_mem_counter[2325] = 4'b0000;
    GSharePlugin_logic_mem_counter[2326] = 4'b0000;
    GSharePlugin_logic_mem_counter[2327] = 4'b0000;
    GSharePlugin_logic_mem_counter[2328] = 4'b0000;
    GSharePlugin_logic_mem_counter[2329] = 4'b0000;
    GSharePlugin_logic_mem_counter[2330] = 4'b0000;
    GSharePlugin_logic_mem_counter[2331] = 4'b0000;
    GSharePlugin_logic_mem_counter[2332] = 4'b0000;
    GSharePlugin_logic_mem_counter[2333] = 4'b0000;
    GSharePlugin_logic_mem_counter[2334] = 4'b0000;
    GSharePlugin_logic_mem_counter[2335] = 4'b0000;
    GSharePlugin_logic_mem_counter[2336] = 4'b0000;
    GSharePlugin_logic_mem_counter[2337] = 4'b0000;
    GSharePlugin_logic_mem_counter[2338] = 4'b0000;
    GSharePlugin_logic_mem_counter[2339] = 4'b0000;
    GSharePlugin_logic_mem_counter[2340] = 4'b0000;
    GSharePlugin_logic_mem_counter[2341] = 4'b0000;
    GSharePlugin_logic_mem_counter[2342] = 4'b0000;
    GSharePlugin_logic_mem_counter[2343] = 4'b0000;
    GSharePlugin_logic_mem_counter[2344] = 4'b0000;
    GSharePlugin_logic_mem_counter[2345] = 4'b0000;
    GSharePlugin_logic_mem_counter[2346] = 4'b0000;
    GSharePlugin_logic_mem_counter[2347] = 4'b0000;
    GSharePlugin_logic_mem_counter[2348] = 4'b0000;
    GSharePlugin_logic_mem_counter[2349] = 4'b0000;
    GSharePlugin_logic_mem_counter[2350] = 4'b0000;
    GSharePlugin_logic_mem_counter[2351] = 4'b0000;
    GSharePlugin_logic_mem_counter[2352] = 4'b0000;
    GSharePlugin_logic_mem_counter[2353] = 4'b0000;
    GSharePlugin_logic_mem_counter[2354] = 4'b0000;
    GSharePlugin_logic_mem_counter[2355] = 4'b0000;
    GSharePlugin_logic_mem_counter[2356] = 4'b0000;
    GSharePlugin_logic_mem_counter[2357] = 4'b0000;
    GSharePlugin_logic_mem_counter[2358] = 4'b0000;
    GSharePlugin_logic_mem_counter[2359] = 4'b0000;
    GSharePlugin_logic_mem_counter[2360] = 4'b0000;
    GSharePlugin_logic_mem_counter[2361] = 4'b0000;
    GSharePlugin_logic_mem_counter[2362] = 4'b0000;
    GSharePlugin_logic_mem_counter[2363] = 4'b0000;
    GSharePlugin_logic_mem_counter[2364] = 4'b0000;
    GSharePlugin_logic_mem_counter[2365] = 4'b0000;
    GSharePlugin_logic_mem_counter[2366] = 4'b0000;
    GSharePlugin_logic_mem_counter[2367] = 4'b0000;
    GSharePlugin_logic_mem_counter[2368] = 4'b0000;
    GSharePlugin_logic_mem_counter[2369] = 4'b0000;
    GSharePlugin_logic_mem_counter[2370] = 4'b0000;
    GSharePlugin_logic_mem_counter[2371] = 4'b0000;
    GSharePlugin_logic_mem_counter[2372] = 4'b0000;
    GSharePlugin_logic_mem_counter[2373] = 4'b0000;
    GSharePlugin_logic_mem_counter[2374] = 4'b0000;
    GSharePlugin_logic_mem_counter[2375] = 4'b0000;
    GSharePlugin_logic_mem_counter[2376] = 4'b0000;
    GSharePlugin_logic_mem_counter[2377] = 4'b0000;
    GSharePlugin_logic_mem_counter[2378] = 4'b0000;
    GSharePlugin_logic_mem_counter[2379] = 4'b0000;
    GSharePlugin_logic_mem_counter[2380] = 4'b0000;
    GSharePlugin_logic_mem_counter[2381] = 4'b0000;
    GSharePlugin_logic_mem_counter[2382] = 4'b0000;
    GSharePlugin_logic_mem_counter[2383] = 4'b0000;
    GSharePlugin_logic_mem_counter[2384] = 4'b0000;
    GSharePlugin_logic_mem_counter[2385] = 4'b0000;
    GSharePlugin_logic_mem_counter[2386] = 4'b0000;
    GSharePlugin_logic_mem_counter[2387] = 4'b0000;
    GSharePlugin_logic_mem_counter[2388] = 4'b0000;
    GSharePlugin_logic_mem_counter[2389] = 4'b0000;
    GSharePlugin_logic_mem_counter[2390] = 4'b0000;
    GSharePlugin_logic_mem_counter[2391] = 4'b0000;
    GSharePlugin_logic_mem_counter[2392] = 4'b0000;
    GSharePlugin_logic_mem_counter[2393] = 4'b0000;
    GSharePlugin_logic_mem_counter[2394] = 4'b0000;
    GSharePlugin_logic_mem_counter[2395] = 4'b0000;
    GSharePlugin_logic_mem_counter[2396] = 4'b0000;
    GSharePlugin_logic_mem_counter[2397] = 4'b0000;
    GSharePlugin_logic_mem_counter[2398] = 4'b0000;
    GSharePlugin_logic_mem_counter[2399] = 4'b0000;
    GSharePlugin_logic_mem_counter[2400] = 4'b0000;
    GSharePlugin_logic_mem_counter[2401] = 4'b0000;
    GSharePlugin_logic_mem_counter[2402] = 4'b0000;
    GSharePlugin_logic_mem_counter[2403] = 4'b0000;
    GSharePlugin_logic_mem_counter[2404] = 4'b0000;
    GSharePlugin_logic_mem_counter[2405] = 4'b0000;
    GSharePlugin_logic_mem_counter[2406] = 4'b0000;
    GSharePlugin_logic_mem_counter[2407] = 4'b0000;
    GSharePlugin_logic_mem_counter[2408] = 4'b0000;
    GSharePlugin_logic_mem_counter[2409] = 4'b0000;
    GSharePlugin_logic_mem_counter[2410] = 4'b0000;
    GSharePlugin_logic_mem_counter[2411] = 4'b0000;
    GSharePlugin_logic_mem_counter[2412] = 4'b0000;
    GSharePlugin_logic_mem_counter[2413] = 4'b0000;
    GSharePlugin_logic_mem_counter[2414] = 4'b0000;
    GSharePlugin_logic_mem_counter[2415] = 4'b0000;
    GSharePlugin_logic_mem_counter[2416] = 4'b0000;
    GSharePlugin_logic_mem_counter[2417] = 4'b0000;
    GSharePlugin_logic_mem_counter[2418] = 4'b0000;
    GSharePlugin_logic_mem_counter[2419] = 4'b0000;
    GSharePlugin_logic_mem_counter[2420] = 4'b0000;
    GSharePlugin_logic_mem_counter[2421] = 4'b0000;
    GSharePlugin_logic_mem_counter[2422] = 4'b0000;
    GSharePlugin_logic_mem_counter[2423] = 4'b0000;
    GSharePlugin_logic_mem_counter[2424] = 4'b0000;
    GSharePlugin_logic_mem_counter[2425] = 4'b0000;
    GSharePlugin_logic_mem_counter[2426] = 4'b0000;
    GSharePlugin_logic_mem_counter[2427] = 4'b0000;
    GSharePlugin_logic_mem_counter[2428] = 4'b0000;
    GSharePlugin_logic_mem_counter[2429] = 4'b0000;
    GSharePlugin_logic_mem_counter[2430] = 4'b0000;
    GSharePlugin_logic_mem_counter[2431] = 4'b0000;
    GSharePlugin_logic_mem_counter[2432] = 4'b0000;
    GSharePlugin_logic_mem_counter[2433] = 4'b0000;
    GSharePlugin_logic_mem_counter[2434] = 4'b0000;
    GSharePlugin_logic_mem_counter[2435] = 4'b0000;
    GSharePlugin_logic_mem_counter[2436] = 4'b0000;
    GSharePlugin_logic_mem_counter[2437] = 4'b0000;
    GSharePlugin_logic_mem_counter[2438] = 4'b0000;
    GSharePlugin_logic_mem_counter[2439] = 4'b0000;
    GSharePlugin_logic_mem_counter[2440] = 4'b0000;
    GSharePlugin_logic_mem_counter[2441] = 4'b0000;
    GSharePlugin_logic_mem_counter[2442] = 4'b0000;
    GSharePlugin_logic_mem_counter[2443] = 4'b0000;
    GSharePlugin_logic_mem_counter[2444] = 4'b0000;
    GSharePlugin_logic_mem_counter[2445] = 4'b0000;
    GSharePlugin_logic_mem_counter[2446] = 4'b0000;
    GSharePlugin_logic_mem_counter[2447] = 4'b0000;
    GSharePlugin_logic_mem_counter[2448] = 4'b0000;
    GSharePlugin_logic_mem_counter[2449] = 4'b0000;
    GSharePlugin_logic_mem_counter[2450] = 4'b0000;
    GSharePlugin_logic_mem_counter[2451] = 4'b0000;
    GSharePlugin_logic_mem_counter[2452] = 4'b0000;
    GSharePlugin_logic_mem_counter[2453] = 4'b0000;
    GSharePlugin_logic_mem_counter[2454] = 4'b0000;
    GSharePlugin_logic_mem_counter[2455] = 4'b0000;
    GSharePlugin_logic_mem_counter[2456] = 4'b0000;
    GSharePlugin_logic_mem_counter[2457] = 4'b0000;
    GSharePlugin_logic_mem_counter[2458] = 4'b0000;
    GSharePlugin_logic_mem_counter[2459] = 4'b0000;
    GSharePlugin_logic_mem_counter[2460] = 4'b0000;
    GSharePlugin_logic_mem_counter[2461] = 4'b0000;
    GSharePlugin_logic_mem_counter[2462] = 4'b0000;
    GSharePlugin_logic_mem_counter[2463] = 4'b0000;
    GSharePlugin_logic_mem_counter[2464] = 4'b0000;
    GSharePlugin_logic_mem_counter[2465] = 4'b0000;
    GSharePlugin_logic_mem_counter[2466] = 4'b0000;
    GSharePlugin_logic_mem_counter[2467] = 4'b0000;
    GSharePlugin_logic_mem_counter[2468] = 4'b0000;
    GSharePlugin_logic_mem_counter[2469] = 4'b0000;
    GSharePlugin_logic_mem_counter[2470] = 4'b0000;
    GSharePlugin_logic_mem_counter[2471] = 4'b0000;
    GSharePlugin_logic_mem_counter[2472] = 4'b0000;
    GSharePlugin_logic_mem_counter[2473] = 4'b0000;
    GSharePlugin_logic_mem_counter[2474] = 4'b0000;
    GSharePlugin_logic_mem_counter[2475] = 4'b0000;
    GSharePlugin_logic_mem_counter[2476] = 4'b0000;
    GSharePlugin_logic_mem_counter[2477] = 4'b0000;
    GSharePlugin_logic_mem_counter[2478] = 4'b0000;
    GSharePlugin_logic_mem_counter[2479] = 4'b0000;
    GSharePlugin_logic_mem_counter[2480] = 4'b0000;
    GSharePlugin_logic_mem_counter[2481] = 4'b0000;
    GSharePlugin_logic_mem_counter[2482] = 4'b0000;
    GSharePlugin_logic_mem_counter[2483] = 4'b0000;
    GSharePlugin_logic_mem_counter[2484] = 4'b0000;
    GSharePlugin_logic_mem_counter[2485] = 4'b0000;
    GSharePlugin_logic_mem_counter[2486] = 4'b0000;
    GSharePlugin_logic_mem_counter[2487] = 4'b0000;
    GSharePlugin_logic_mem_counter[2488] = 4'b0000;
    GSharePlugin_logic_mem_counter[2489] = 4'b0000;
    GSharePlugin_logic_mem_counter[2490] = 4'b0000;
    GSharePlugin_logic_mem_counter[2491] = 4'b0000;
    GSharePlugin_logic_mem_counter[2492] = 4'b0000;
    GSharePlugin_logic_mem_counter[2493] = 4'b0000;
    GSharePlugin_logic_mem_counter[2494] = 4'b0000;
    GSharePlugin_logic_mem_counter[2495] = 4'b0000;
    GSharePlugin_logic_mem_counter[2496] = 4'b0000;
    GSharePlugin_logic_mem_counter[2497] = 4'b0000;
    GSharePlugin_logic_mem_counter[2498] = 4'b0000;
    GSharePlugin_logic_mem_counter[2499] = 4'b0000;
    GSharePlugin_logic_mem_counter[2500] = 4'b0000;
    GSharePlugin_logic_mem_counter[2501] = 4'b0000;
    GSharePlugin_logic_mem_counter[2502] = 4'b0000;
    GSharePlugin_logic_mem_counter[2503] = 4'b0000;
    GSharePlugin_logic_mem_counter[2504] = 4'b0000;
    GSharePlugin_logic_mem_counter[2505] = 4'b0000;
    GSharePlugin_logic_mem_counter[2506] = 4'b0000;
    GSharePlugin_logic_mem_counter[2507] = 4'b0000;
    GSharePlugin_logic_mem_counter[2508] = 4'b0000;
    GSharePlugin_logic_mem_counter[2509] = 4'b0000;
    GSharePlugin_logic_mem_counter[2510] = 4'b0000;
    GSharePlugin_logic_mem_counter[2511] = 4'b0000;
    GSharePlugin_logic_mem_counter[2512] = 4'b0000;
    GSharePlugin_logic_mem_counter[2513] = 4'b0000;
    GSharePlugin_logic_mem_counter[2514] = 4'b0000;
    GSharePlugin_logic_mem_counter[2515] = 4'b0000;
    GSharePlugin_logic_mem_counter[2516] = 4'b0000;
    GSharePlugin_logic_mem_counter[2517] = 4'b0000;
    GSharePlugin_logic_mem_counter[2518] = 4'b0000;
    GSharePlugin_logic_mem_counter[2519] = 4'b0000;
    GSharePlugin_logic_mem_counter[2520] = 4'b0000;
    GSharePlugin_logic_mem_counter[2521] = 4'b0000;
    GSharePlugin_logic_mem_counter[2522] = 4'b0000;
    GSharePlugin_logic_mem_counter[2523] = 4'b0000;
    GSharePlugin_logic_mem_counter[2524] = 4'b0000;
    GSharePlugin_logic_mem_counter[2525] = 4'b0000;
    GSharePlugin_logic_mem_counter[2526] = 4'b0000;
    GSharePlugin_logic_mem_counter[2527] = 4'b0000;
    GSharePlugin_logic_mem_counter[2528] = 4'b0000;
    GSharePlugin_logic_mem_counter[2529] = 4'b0000;
    GSharePlugin_logic_mem_counter[2530] = 4'b0000;
    GSharePlugin_logic_mem_counter[2531] = 4'b0000;
    GSharePlugin_logic_mem_counter[2532] = 4'b0000;
    GSharePlugin_logic_mem_counter[2533] = 4'b0000;
    GSharePlugin_logic_mem_counter[2534] = 4'b0000;
    GSharePlugin_logic_mem_counter[2535] = 4'b0000;
    GSharePlugin_logic_mem_counter[2536] = 4'b0000;
    GSharePlugin_logic_mem_counter[2537] = 4'b0000;
    GSharePlugin_logic_mem_counter[2538] = 4'b0000;
    GSharePlugin_logic_mem_counter[2539] = 4'b0000;
    GSharePlugin_logic_mem_counter[2540] = 4'b0000;
    GSharePlugin_logic_mem_counter[2541] = 4'b0000;
    GSharePlugin_logic_mem_counter[2542] = 4'b0000;
    GSharePlugin_logic_mem_counter[2543] = 4'b0000;
    GSharePlugin_logic_mem_counter[2544] = 4'b0000;
    GSharePlugin_logic_mem_counter[2545] = 4'b0000;
    GSharePlugin_logic_mem_counter[2546] = 4'b0000;
    GSharePlugin_logic_mem_counter[2547] = 4'b0000;
    GSharePlugin_logic_mem_counter[2548] = 4'b0000;
    GSharePlugin_logic_mem_counter[2549] = 4'b0000;
    GSharePlugin_logic_mem_counter[2550] = 4'b0000;
    GSharePlugin_logic_mem_counter[2551] = 4'b0000;
    GSharePlugin_logic_mem_counter[2552] = 4'b0000;
    GSharePlugin_logic_mem_counter[2553] = 4'b0000;
    GSharePlugin_logic_mem_counter[2554] = 4'b0000;
    GSharePlugin_logic_mem_counter[2555] = 4'b0000;
    GSharePlugin_logic_mem_counter[2556] = 4'b0000;
    GSharePlugin_logic_mem_counter[2557] = 4'b0000;
    GSharePlugin_logic_mem_counter[2558] = 4'b0000;
    GSharePlugin_logic_mem_counter[2559] = 4'b0000;
    GSharePlugin_logic_mem_counter[2560] = 4'b0000;
    GSharePlugin_logic_mem_counter[2561] = 4'b0000;
    GSharePlugin_logic_mem_counter[2562] = 4'b0000;
    GSharePlugin_logic_mem_counter[2563] = 4'b0000;
    GSharePlugin_logic_mem_counter[2564] = 4'b0000;
    GSharePlugin_logic_mem_counter[2565] = 4'b0000;
    GSharePlugin_logic_mem_counter[2566] = 4'b0000;
    GSharePlugin_logic_mem_counter[2567] = 4'b0000;
    GSharePlugin_logic_mem_counter[2568] = 4'b0000;
    GSharePlugin_logic_mem_counter[2569] = 4'b0000;
    GSharePlugin_logic_mem_counter[2570] = 4'b0000;
    GSharePlugin_logic_mem_counter[2571] = 4'b0000;
    GSharePlugin_logic_mem_counter[2572] = 4'b0000;
    GSharePlugin_logic_mem_counter[2573] = 4'b0000;
    GSharePlugin_logic_mem_counter[2574] = 4'b0000;
    GSharePlugin_logic_mem_counter[2575] = 4'b0000;
    GSharePlugin_logic_mem_counter[2576] = 4'b0000;
    GSharePlugin_logic_mem_counter[2577] = 4'b0000;
    GSharePlugin_logic_mem_counter[2578] = 4'b0000;
    GSharePlugin_logic_mem_counter[2579] = 4'b0000;
    GSharePlugin_logic_mem_counter[2580] = 4'b0000;
    GSharePlugin_logic_mem_counter[2581] = 4'b0000;
    GSharePlugin_logic_mem_counter[2582] = 4'b0000;
    GSharePlugin_logic_mem_counter[2583] = 4'b0000;
    GSharePlugin_logic_mem_counter[2584] = 4'b0000;
    GSharePlugin_logic_mem_counter[2585] = 4'b0000;
    GSharePlugin_logic_mem_counter[2586] = 4'b0000;
    GSharePlugin_logic_mem_counter[2587] = 4'b0000;
    GSharePlugin_logic_mem_counter[2588] = 4'b0000;
    GSharePlugin_logic_mem_counter[2589] = 4'b0000;
    GSharePlugin_logic_mem_counter[2590] = 4'b0000;
    GSharePlugin_logic_mem_counter[2591] = 4'b0000;
    GSharePlugin_logic_mem_counter[2592] = 4'b0000;
    GSharePlugin_logic_mem_counter[2593] = 4'b0000;
    GSharePlugin_logic_mem_counter[2594] = 4'b0000;
    GSharePlugin_logic_mem_counter[2595] = 4'b0000;
    GSharePlugin_logic_mem_counter[2596] = 4'b0000;
    GSharePlugin_logic_mem_counter[2597] = 4'b0000;
    GSharePlugin_logic_mem_counter[2598] = 4'b0000;
    GSharePlugin_logic_mem_counter[2599] = 4'b0000;
    GSharePlugin_logic_mem_counter[2600] = 4'b0000;
    GSharePlugin_logic_mem_counter[2601] = 4'b0000;
    GSharePlugin_logic_mem_counter[2602] = 4'b0000;
    GSharePlugin_logic_mem_counter[2603] = 4'b0000;
    GSharePlugin_logic_mem_counter[2604] = 4'b0000;
    GSharePlugin_logic_mem_counter[2605] = 4'b0000;
    GSharePlugin_logic_mem_counter[2606] = 4'b0000;
    GSharePlugin_logic_mem_counter[2607] = 4'b0000;
    GSharePlugin_logic_mem_counter[2608] = 4'b0000;
    GSharePlugin_logic_mem_counter[2609] = 4'b0000;
    GSharePlugin_logic_mem_counter[2610] = 4'b0000;
    GSharePlugin_logic_mem_counter[2611] = 4'b0000;
    GSharePlugin_logic_mem_counter[2612] = 4'b0000;
    GSharePlugin_logic_mem_counter[2613] = 4'b0000;
    GSharePlugin_logic_mem_counter[2614] = 4'b0000;
    GSharePlugin_logic_mem_counter[2615] = 4'b0000;
    GSharePlugin_logic_mem_counter[2616] = 4'b0000;
    GSharePlugin_logic_mem_counter[2617] = 4'b0000;
    GSharePlugin_logic_mem_counter[2618] = 4'b0000;
    GSharePlugin_logic_mem_counter[2619] = 4'b0000;
    GSharePlugin_logic_mem_counter[2620] = 4'b0000;
    GSharePlugin_logic_mem_counter[2621] = 4'b0000;
    GSharePlugin_logic_mem_counter[2622] = 4'b0000;
    GSharePlugin_logic_mem_counter[2623] = 4'b0000;
    GSharePlugin_logic_mem_counter[2624] = 4'b0000;
    GSharePlugin_logic_mem_counter[2625] = 4'b0000;
    GSharePlugin_logic_mem_counter[2626] = 4'b0000;
    GSharePlugin_logic_mem_counter[2627] = 4'b0000;
    GSharePlugin_logic_mem_counter[2628] = 4'b0000;
    GSharePlugin_logic_mem_counter[2629] = 4'b0000;
    GSharePlugin_logic_mem_counter[2630] = 4'b0000;
    GSharePlugin_logic_mem_counter[2631] = 4'b0000;
    GSharePlugin_logic_mem_counter[2632] = 4'b0000;
    GSharePlugin_logic_mem_counter[2633] = 4'b0000;
    GSharePlugin_logic_mem_counter[2634] = 4'b0000;
    GSharePlugin_logic_mem_counter[2635] = 4'b0000;
    GSharePlugin_logic_mem_counter[2636] = 4'b0000;
    GSharePlugin_logic_mem_counter[2637] = 4'b0000;
    GSharePlugin_logic_mem_counter[2638] = 4'b0000;
    GSharePlugin_logic_mem_counter[2639] = 4'b0000;
    GSharePlugin_logic_mem_counter[2640] = 4'b0000;
    GSharePlugin_logic_mem_counter[2641] = 4'b0000;
    GSharePlugin_logic_mem_counter[2642] = 4'b0000;
    GSharePlugin_logic_mem_counter[2643] = 4'b0000;
    GSharePlugin_logic_mem_counter[2644] = 4'b0000;
    GSharePlugin_logic_mem_counter[2645] = 4'b0000;
    GSharePlugin_logic_mem_counter[2646] = 4'b0000;
    GSharePlugin_logic_mem_counter[2647] = 4'b0000;
    GSharePlugin_logic_mem_counter[2648] = 4'b0000;
    GSharePlugin_logic_mem_counter[2649] = 4'b0000;
    GSharePlugin_logic_mem_counter[2650] = 4'b0000;
    GSharePlugin_logic_mem_counter[2651] = 4'b0000;
    GSharePlugin_logic_mem_counter[2652] = 4'b0000;
    GSharePlugin_logic_mem_counter[2653] = 4'b0000;
    GSharePlugin_logic_mem_counter[2654] = 4'b0000;
    GSharePlugin_logic_mem_counter[2655] = 4'b0000;
    GSharePlugin_logic_mem_counter[2656] = 4'b0000;
    GSharePlugin_logic_mem_counter[2657] = 4'b0000;
    GSharePlugin_logic_mem_counter[2658] = 4'b0000;
    GSharePlugin_logic_mem_counter[2659] = 4'b0000;
    GSharePlugin_logic_mem_counter[2660] = 4'b0000;
    GSharePlugin_logic_mem_counter[2661] = 4'b0000;
    GSharePlugin_logic_mem_counter[2662] = 4'b0000;
    GSharePlugin_logic_mem_counter[2663] = 4'b0000;
    GSharePlugin_logic_mem_counter[2664] = 4'b0000;
    GSharePlugin_logic_mem_counter[2665] = 4'b0000;
    GSharePlugin_logic_mem_counter[2666] = 4'b0000;
    GSharePlugin_logic_mem_counter[2667] = 4'b0000;
    GSharePlugin_logic_mem_counter[2668] = 4'b0000;
    GSharePlugin_logic_mem_counter[2669] = 4'b0000;
    GSharePlugin_logic_mem_counter[2670] = 4'b0000;
    GSharePlugin_logic_mem_counter[2671] = 4'b0000;
    GSharePlugin_logic_mem_counter[2672] = 4'b0000;
    GSharePlugin_logic_mem_counter[2673] = 4'b0000;
    GSharePlugin_logic_mem_counter[2674] = 4'b0000;
    GSharePlugin_logic_mem_counter[2675] = 4'b0000;
    GSharePlugin_logic_mem_counter[2676] = 4'b0000;
    GSharePlugin_logic_mem_counter[2677] = 4'b0000;
    GSharePlugin_logic_mem_counter[2678] = 4'b0000;
    GSharePlugin_logic_mem_counter[2679] = 4'b0000;
    GSharePlugin_logic_mem_counter[2680] = 4'b0000;
    GSharePlugin_logic_mem_counter[2681] = 4'b0000;
    GSharePlugin_logic_mem_counter[2682] = 4'b0000;
    GSharePlugin_logic_mem_counter[2683] = 4'b0000;
    GSharePlugin_logic_mem_counter[2684] = 4'b0000;
    GSharePlugin_logic_mem_counter[2685] = 4'b0000;
    GSharePlugin_logic_mem_counter[2686] = 4'b0000;
    GSharePlugin_logic_mem_counter[2687] = 4'b0000;
    GSharePlugin_logic_mem_counter[2688] = 4'b0000;
    GSharePlugin_logic_mem_counter[2689] = 4'b0000;
    GSharePlugin_logic_mem_counter[2690] = 4'b0000;
    GSharePlugin_logic_mem_counter[2691] = 4'b0000;
    GSharePlugin_logic_mem_counter[2692] = 4'b0000;
    GSharePlugin_logic_mem_counter[2693] = 4'b0000;
    GSharePlugin_logic_mem_counter[2694] = 4'b0000;
    GSharePlugin_logic_mem_counter[2695] = 4'b0000;
    GSharePlugin_logic_mem_counter[2696] = 4'b0000;
    GSharePlugin_logic_mem_counter[2697] = 4'b0000;
    GSharePlugin_logic_mem_counter[2698] = 4'b0000;
    GSharePlugin_logic_mem_counter[2699] = 4'b0000;
    GSharePlugin_logic_mem_counter[2700] = 4'b0000;
    GSharePlugin_logic_mem_counter[2701] = 4'b0000;
    GSharePlugin_logic_mem_counter[2702] = 4'b0000;
    GSharePlugin_logic_mem_counter[2703] = 4'b0000;
    GSharePlugin_logic_mem_counter[2704] = 4'b0000;
    GSharePlugin_logic_mem_counter[2705] = 4'b0000;
    GSharePlugin_logic_mem_counter[2706] = 4'b0000;
    GSharePlugin_logic_mem_counter[2707] = 4'b0000;
    GSharePlugin_logic_mem_counter[2708] = 4'b0000;
    GSharePlugin_logic_mem_counter[2709] = 4'b0000;
    GSharePlugin_logic_mem_counter[2710] = 4'b0000;
    GSharePlugin_logic_mem_counter[2711] = 4'b0000;
    GSharePlugin_logic_mem_counter[2712] = 4'b0000;
    GSharePlugin_logic_mem_counter[2713] = 4'b0000;
    GSharePlugin_logic_mem_counter[2714] = 4'b0000;
    GSharePlugin_logic_mem_counter[2715] = 4'b0000;
    GSharePlugin_logic_mem_counter[2716] = 4'b0000;
    GSharePlugin_logic_mem_counter[2717] = 4'b0000;
    GSharePlugin_logic_mem_counter[2718] = 4'b0000;
    GSharePlugin_logic_mem_counter[2719] = 4'b0000;
    GSharePlugin_logic_mem_counter[2720] = 4'b0000;
    GSharePlugin_logic_mem_counter[2721] = 4'b0000;
    GSharePlugin_logic_mem_counter[2722] = 4'b0000;
    GSharePlugin_logic_mem_counter[2723] = 4'b0000;
    GSharePlugin_logic_mem_counter[2724] = 4'b0000;
    GSharePlugin_logic_mem_counter[2725] = 4'b0000;
    GSharePlugin_logic_mem_counter[2726] = 4'b0000;
    GSharePlugin_logic_mem_counter[2727] = 4'b0000;
    GSharePlugin_logic_mem_counter[2728] = 4'b0000;
    GSharePlugin_logic_mem_counter[2729] = 4'b0000;
    GSharePlugin_logic_mem_counter[2730] = 4'b0000;
    GSharePlugin_logic_mem_counter[2731] = 4'b0000;
    GSharePlugin_logic_mem_counter[2732] = 4'b0000;
    GSharePlugin_logic_mem_counter[2733] = 4'b0000;
    GSharePlugin_logic_mem_counter[2734] = 4'b0000;
    GSharePlugin_logic_mem_counter[2735] = 4'b0000;
    GSharePlugin_logic_mem_counter[2736] = 4'b0000;
    GSharePlugin_logic_mem_counter[2737] = 4'b0000;
    GSharePlugin_logic_mem_counter[2738] = 4'b0000;
    GSharePlugin_logic_mem_counter[2739] = 4'b0000;
    GSharePlugin_logic_mem_counter[2740] = 4'b0000;
    GSharePlugin_logic_mem_counter[2741] = 4'b0000;
    GSharePlugin_logic_mem_counter[2742] = 4'b0000;
    GSharePlugin_logic_mem_counter[2743] = 4'b0000;
    GSharePlugin_logic_mem_counter[2744] = 4'b0000;
    GSharePlugin_logic_mem_counter[2745] = 4'b0000;
    GSharePlugin_logic_mem_counter[2746] = 4'b0000;
    GSharePlugin_logic_mem_counter[2747] = 4'b0000;
    GSharePlugin_logic_mem_counter[2748] = 4'b0000;
    GSharePlugin_logic_mem_counter[2749] = 4'b0000;
    GSharePlugin_logic_mem_counter[2750] = 4'b0000;
    GSharePlugin_logic_mem_counter[2751] = 4'b0000;
    GSharePlugin_logic_mem_counter[2752] = 4'b0000;
    GSharePlugin_logic_mem_counter[2753] = 4'b0000;
    GSharePlugin_logic_mem_counter[2754] = 4'b0000;
    GSharePlugin_logic_mem_counter[2755] = 4'b0000;
    GSharePlugin_logic_mem_counter[2756] = 4'b0000;
    GSharePlugin_logic_mem_counter[2757] = 4'b0000;
    GSharePlugin_logic_mem_counter[2758] = 4'b0000;
    GSharePlugin_logic_mem_counter[2759] = 4'b0000;
    GSharePlugin_logic_mem_counter[2760] = 4'b0000;
    GSharePlugin_logic_mem_counter[2761] = 4'b0000;
    GSharePlugin_logic_mem_counter[2762] = 4'b0000;
    GSharePlugin_logic_mem_counter[2763] = 4'b0000;
    GSharePlugin_logic_mem_counter[2764] = 4'b0000;
    GSharePlugin_logic_mem_counter[2765] = 4'b0000;
    GSharePlugin_logic_mem_counter[2766] = 4'b0000;
    GSharePlugin_logic_mem_counter[2767] = 4'b0000;
    GSharePlugin_logic_mem_counter[2768] = 4'b0000;
    GSharePlugin_logic_mem_counter[2769] = 4'b0000;
    GSharePlugin_logic_mem_counter[2770] = 4'b0000;
    GSharePlugin_logic_mem_counter[2771] = 4'b0000;
    GSharePlugin_logic_mem_counter[2772] = 4'b0000;
    GSharePlugin_logic_mem_counter[2773] = 4'b0000;
    GSharePlugin_logic_mem_counter[2774] = 4'b0000;
    GSharePlugin_logic_mem_counter[2775] = 4'b0000;
    GSharePlugin_logic_mem_counter[2776] = 4'b0000;
    GSharePlugin_logic_mem_counter[2777] = 4'b0000;
    GSharePlugin_logic_mem_counter[2778] = 4'b0000;
    GSharePlugin_logic_mem_counter[2779] = 4'b0000;
    GSharePlugin_logic_mem_counter[2780] = 4'b0000;
    GSharePlugin_logic_mem_counter[2781] = 4'b0000;
    GSharePlugin_logic_mem_counter[2782] = 4'b0000;
    GSharePlugin_logic_mem_counter[2783] = 4'b0000;
    GSharePlugin_logic_mem_counter[2784] = 4'b0000;
    GSharePlugin_logic_mem_counter[2785] = 4'b0000;
    GSharePlugin_logic_mem_counter[2786] = 4'b0000;
    GSharePlugin_logic_mem_counter[2787] = 4'b0000;
    GSharePlugin_logic_mem_counter[2788] = 4'b0000;
    GSharePlugin_logic_mem_counter[2789] = 4'b0000;
    GSharePlugin_logic_mem_counter[2790] = 4'b0000;
    GSharePlugin_logic_mem_counter[2791] = 4'b0000;
    GSharePlugin_logic_mem_counter[2792] = 4'b0000;
    GSharePlugin_logic_mem_counter[2793] = 4'b0000;
    GSharePlugin_logic_mem_counter[2794] = 4'b0000;
    GSharePlugin_logic_mem_counter[2795] = 4'b0000;
    GSharePlugin_logic_mem_counter[2796] = 4'b0000;
    GSharePlugin_logic_mem_counter[2797] = 4'b0000;
    GSharePlugin_logic_mem_counter[2798] = 4'b0000;
    GSharePlugin_logic_mem_counter[2799] = 4'b0000;
    GSharePlugin_logic_mem_counter[2800] = 4'b0000;
    GSharePlugin_logic_mem_counter[2801] = 4'b0000;
    GSharePlugin_logic_mem_counter[2802] = 4'b0000;
    GSharePlugin_logic_mem_counter[2803] = 4'b0000;
    GSharePlugin_logic_mem_counter[2804] = 4'b0000;
    GSharePlugin_logic_mem_counter[2805] = 4'b0000;
    GSharePlugin_logic_mem_counter[2806] = 4'b0000;
    GSharePlugin_logic_mem_counter[2807] = 4'b0000;
    GSharePlugin_logic_mem_counter[2808] = 4'b0000;
    GSharePlugin_logic_mem_counter[2809] = 4'b0000;
    GSharePlugin_logic_mem_counter[2810] = 4'b0000;
    GSharePlugin_logic_mem_counter[2811] = 4'b0000;
    GSharePlugin_logic_mem_counter[2812] = 4'b0000;
    GSharePlugin_logic_mem_counter[2813] = 4'b0000;
    GSharePlugin_logic_mem_counter[2814] = 4'b0000;
    GSharePlugin_logic_mem_counter[2815] = 4'b0000;
    GSharePlugin_logic_mem_counter[2816] = 4'b0000;
    GSharePlugin_logic_mem_counter[2817] = 4'b0000;
    GSharePlugin_logic_mem_counter[2818] = 4'b0000;
    GSharePlugin_logic_mem_counter[2819] = 4'b0000;
    GSharePlugin_logic_mem_counter[2820] = 4'b0000;
    GSharePlugin_logic_mem_counter[2821] = 4'b0000;
    GSharePlugin_logic_mem_counter[2822] = 4'b0000;
    GSharePlugin_logic_mem_counter[2823] = 4'b0000;
    GSharePlugin_logic_mem_counter[2824] = 4'b0000;
    GSharePlugin_logic_mem_counter[2825] = 4'b0000;
    GSharePlugin_logic_mem_counter[2826] = 4'b0000;
    GSharePlugin_logic_mem_counter[2827] = 4'b0000;
    GSharePlugin_logic_mem_counter[2828] = 4'b0000;
    GSharePlugin_logic_mem_counter[2829] = 4'b0000;
    GSharePlugin_logic_mem_counter[2830] = 4'b0000;
    GSharePlugin_logic_mem_counter[2831] = 4'b0000;
    GSharePlugin_logic_mem_counter[2832] = 4'b0000;
    GSharePlugin_logic_mem_counter[2833] = 4'b0000;
    GSharePlugin_logic_mem_counter[2834] = 4'b0000;
    GSharePlugin_logic_mem_counter[2835] = 4'b0000;
    GSharePlugin_logic_mem_counter[2836] = 4'b0000;
    GSharePlugin_logic_mem_counter[2837] = 4'b0000;
    GSharePlugin_logic_mem_counter[2838] = 4'b0000;
    GSharePlugin_logic_mem_counter[2839] = 4'b0000;
    GSharePlugin_logic_mem_counter[2840] = 4'b0000;
    GSharePlugin_logic_mem_counter[2841] = 4'b0000;
    GSharePlugin_logic_mem_counter[2842] = 4'b0000;
    GSharePlugin_logic_mem_counter[2843] = 4'b0000;
    GSharePlugin_logic_mem_counter[2844] = 4'b0000;
    GSharePlugin_logic_mem_counter[2845] = 4'b0000;
    GSharePlugin_logic_mem_counter[2846] = 4'b0000;
    GSharePlugin_logic_mem_counter[2847] = 4'b0000;
    GSharePlugin_logic_mem_counter[2848] = 4'b0000;
    GSharePlugin_logic_mem_counter[2849] = 4'b0000;
    GSharePlugin_logic_mem_counter[2850] = 4'b0000;
    GSharePlugin_logic_mem_counter[2851] = 4'b0000;
    GSharePlugin_logic_mem_counter[2852] = 4'b0000;
    GSharePlugin_logic_mem_counter[2853] = 4'b0000;
    GSharePlugin_logic_mem_counter[2854] = 4'b0000;
    GSharePlugin_logic_mem_counter[2855] = 4'b0000;
    GSharePlugin_logic_mem_counter[2856] = 4'b0000;
    GSharePlugin_logic_mem_counter[2857] = 4'b0000;
    GSharePlugin_logic_mem_counter[2858] = 4'b0000;
    GSharePlugin_logic_mem_counter[2859] = 4'b0000;
    GSharePlugin_logic_mem_counter[2860] = 4'b0000;
    GSharePlugin_logic_mem_counter[2861] = 4'b0000;
    GSharePlugin_logic_mem_counter[2862] = 4'b0000;
    GSharePlugin_logic_mem_counter[2863] = 4'b0000;
    GSharePlugin_logic_mem_counter[2864] = 4'b0000;
    GSharePlugin_logic_mem_counter[2865] = 4'b0000;
    GSharePlugin_logic_mem_counter[2866] = 4'b0000;
    GSharePlugin_logic_mem_counter[2867] = 4'b0000;
    GSharePlugin_logic_mem_counter[2868] = 4'b0000;
    GSharePlugin_logic_mem_counter[2869] = 4'b0000;
    GSharePlugin_logic_mem_counter[2870] = 4'b0000;
    GSharePlugin_logic_mem_counter[2871] = 4'b0000;
    GSharePlugin_logic_mem_counter[2872] = 4'b0000;
    GSharePlugin_logic_mem_counter[2873] = 4'b0000;
    GSharePlugin_logic_mem_counter[2874] = 4'b0000;
    GSharePlugin_logic_mem_counter[2875] = 4'b0000;
    GSharePlugin_logic_mem_counter[2876] = 4'b0000;
    GSharePlugin_logic_mem_counter[2877] = 4'b0000;
    GSharePlugin_logic_mem_counter[2878] = 4'b0000;
    GSharePlugin_logic_mem_counter[2879] = 4'b0000;
    GSharePlugin_logic_mem_counter[2880] = 4'b0000;
    GSharePlugin_logic_mem_counter[2881] = 4'b0000;
    GSharePlugin_logic_mem_counter[2882] = 4'b0000;
    GSharePlugin_logic_mem_counter[2883] = 4'b0000;
    GSharePlugin_logic_mem_counter[2884] = 4'b0000;
    GSharePlugin_logic_mem_counter[2885] = 4'b0000;
    GSharePlugin_logic_mem_counter[2886] = 4'b0000;
    GSharePlugin_logic_mem_counter[2887] = 4'b0000;
    GSharePlugin_logic_mem_counter[2888] = 4'b0000;
    GSharePlugin_logic_mem_counter[2889] = 4'b0000;
    GSharePlugin_logic_mem_counter[2890] = 4'b0000;
    GSharePlugin_logic_mem_counter[2891] = 4'b0000;
    GSharePlugin_logic_mem_counter[2892] = 4'b0000;
    GSharePlugin_logic_mem_counter[2893] = 4'b0000;
    GSharePlugin_logic_mem_counter[2894] = 4'b0000;
    GSharePlugin_logic_mem_counter[2895] = 4'b0000;
    GSharePlugin_logic_mem_counter[2896] = 4'b0000;
    GSharePlugin_logic_mem_counter[2897] = 4'b0000;
    GSharePlugin_logic_mem_counter[2898] = 4'b0000;
    GSharePlugin_logic_mem_counter[2899] = 4'b0000;
    GSharePlugin_logic_mem_counter[2900] = 4'b0000;
    GSharePlugin_logic_mem_counter[2901] = 4'b0000;
    GSharePlugin_logic_mem_counter[2902] = 4'b0000;
    GSharePlugin_logic_mem_counter[2903] = 4'b0000;
    GSharePlugin_logic_mem_counter[2904] = 4'b0000;
    GSharePlugin_logic_mem_counter[2905] = 4'b0000;
    GSharePlugin_logic_mem_counter[2906] = 4'b0000;
    GSharePlugin_logic_mem_counter[2907] = 4'b0000;
    GSharePlugin_logic_mem_counter[2908] = 4'b0000;
    GSharePlugin_logic_mem_counter[2909] = 4'b0000;
    GSharePlugin_logic_mem_counter[2910] = 4'b0000;
    GSharePlugin_logic_mem_counter[2911] = 4'b0000;
    GSharePlugin_logic_mem_counter[2912] = 4'b0000;
    GSharePlugin_logic_mem_counter[2913] = 4'b0000;
    GSharePlugin_logic_mem_counter[2914] = 4'b0000;
    GSharePlugin_logic_mem_counter[2915] = 4'b0000;
    GSharePlugin_logic_mem_counter[2916] = 4'b0000;
    GSharePlugin_logic_mem_counter[2917] = 4'b0000;
    GSharePlugin_logic_mem_counter[2918] = 4'b0000;
    GSharePlugin_logic_mem_counter[2919] = 4'b0000;
    GSharePlugin_logic_mem_counter[2920] = 4'b0000;
    GSharePlugin_logic_mem_counter[2921] = 4'b0000;
    GSharePlugin_logic_mem_counter[2922] = 4'b0000;
    GSharePlugin_logic_mem_counter[2923] = 4'b0000;
    GSharePlugin_logic_mem_counter[2924] = 4'b0000;
    GSharePlugin_logic_mem_counter[2925] = 4'b0000;
    GSharePlugin_logic_mem_counter[2926] = 4'b0000;
    GSharePlugin_logic_mem_counter[2927] = 4'b0000;
    GSharePlugin_logic_mem_counter[2928] = 4'b0000;
    GSharePlugin_logic_mem_counter[2929] = 4'b0000;
    GSharePlugin_logic_mem_counter[2930] = 4'b0000;
    GSharePlugin_logic_mem_counter[2931] = 4'b0000;
    GSharePlugin_logic_mem_counter[2932] = 4'b0000;
    GSharePlugin_logic_mem_counter[2933] = 4'b0000;
    GSharePlugin_logic_mem_counter[2934] = 4'b0000;
    GSharePlugin_logic_mem_counter[2935] = 4'b0000;
    GSharePlugin_logic_mem_counter[2936] = 4'b0000;
    GSharePlugin_logic_mem_counter[2937] = 4'b0000;
    GSharePlugin_logic_mem_counter[2938] = 4'b0000;
    GSharePlugin_logic_mem_counter[2939] = 4'b0000;
    GSharePlugin_logic_mem_counter[2940] = 4'b0000;
    GSharePlugin_logic_mem_counter[2941] = 4'b0000;
    GSharePlugin_logic_mem_counter[2942] = 4'b0000;
    GSharePlugin_logic_mem_counter[2943] = 4'b0000;
    GSharePlugin_logic_mem_counter[2944] = 4'b0000;
    GSharePlugin_logic_mem_counter[2945] = 4'b0000;
    GSharePlugin_logic_mem_counter[2946] = 4'b0000;
    GSharePlugin_logic_mem_counter[2947] = 4'b0000;
    GSharePlugin_logic_mem_counter[2948] = 4'b0000;
    GSharePlugin_logic_mem_counter[2949] = 4'b0000;
    GSharePlugin_logic_mem_counter[2950] = 4'b0000;
    GSharePlugin_logic_mem_counter[2951] = 4'b0000;
    GSharePlugin_logic_mem_counter[2952] = 4'b0000;
    GSharePlugin_logic_mem_counter[2953] = 4'b0000;
    GSharePlugin_logic_mem_counter[2954] = 4'b0000;
    GSharePlugin_logic_mem_counter[2955] = 4'b0000;
    GSharePlugin_logic_mem_counter[2956] = 4'b0000;
    GSharePlugin_logic_mem_counter[2957] = 4'b0000;
    GSharePlugin_logic_mem_counter[2958] = 4'b0000;
    GSharePlugin_logic_mem_counter[2959] = 4'b0000;
    GSharePlugin_logic_mem_counter[2960] = 4'b0000;
    GSharePlugin_logic_mem_counter[2961] = 4'b0000;
    GSharePlugin_logic_mem_counter[2962] = 4'b0000;
    GSharePlugin_logic_mem_counter[2963] = 4'b0000;
    GSharePlugin_logic_mem_counter[2964] = 4'b0000;
    GSharePlugin_logic_mem_counter[2965] = 4'b0000;
    GSharePlugin_logic_mem_counter[2966] = 4'b0000;
    GSharePlugin_logic_mem_counter[2967] = 4'b0000;
    GSharePlugin_logic_mem_counter[2968] = 4'b0000;
    GSharePlugin_logic_mem_counter[2969] = 4'b0000;
    GSharePlugin_logic_mem_counter[2970] = 4'b0000;
    GSharePlugin_logic_mem_counter[2971] = 4'b0000;
    GSharePlugin_logic_mem_counter[2972] = 4'b0000;
    GSharePlugin_logic_mem_counter[2973] = 4'b0000;
    GSharePlugin_logic_mem_counter[2974] = 4'b0000;
    GSharePlugin_logic_mem_counter[2975] = 4'b0000;
    GSharePlugin_logic_mem_counter[2976] = 4'b0000;
    GSharePlugin_logic_mem_counter[2977] = 4'b0000;
    GSharePlugin_logic_mem_counter[2978] = 4'b0000;
    GSharePlugin_logic_mem_counter[2979] = 4'b0000;
    GSharePlugin_logic_mem_counter[2980] = 4'b0000;
    GSharePlugin_logic_mem_counter[2981] = 4'b0000;
    GSharePlugin_logic_mem_counter[2982] = 4'b0000;
    GSharePlugin_logic_mem_counter[2983] = 4'b0000;
    GSharePlugin_logic_mem_counter[2984] = 4'b0000;
    GSharePlugin_logic_mem_counter[2985] = 4'b0000;
    GSharePlugin_logic_mem_counter[2986] = 4'b0000;
    GSharePlugin_logic_mem_counter[2987] = 4'b0000;
    GSharePlugin_logic_mem_counter[2988] = 4'b0000;
    GSharePlugin_logic_mem_counter[2989] = 4'b0000;
    GSharePlugin_logic_mem_counter[2990] = 4'b0000;
    GSharePlugin_logic_mem_counter[2991] = 4'b0000;
    GSharePlugin_logic_mem_counter[2992] = 4'b0000;
    GSharePlugin_logic_mem_counter[2993] = 4'b0000;
    GSharePlugin_logic_mem_counter[2994] = 4'b0000;
    GSharePlugin_logic_mem_counter[2995] = 4'b0000;
    GSharePlugin_logic_mem_counter[2996] = 4'b0000;
    GSharePlugin_logic_mem_counter[2997] = 4'b0000;
    GSharePlugin_logic_mem_counter[2998] = 4'b0000;
    GSharePlugin_logic_mem_counter[2999] = 4'b0000;
    GSharePlugin_logic_mem_counter[3000] = 4'b0000;
    GSharePlugin_logic_mem_counter[3001] = 4'b0000;
    GSharePlugin_logic_mem_counter[3002] = 4'b0000;
    GSharePlugin_logic_mem_counter[3003] = 4'b0000;
    GSharePlugin_logic_mem_counter[3004] = 4'b0000;
    GSharePlugin_logic_mem_counter[3005] = 4'b0000;
    GSharePlugin_logic_mem_counter[3006] = 4'b0000;
    GSharePlugin_logic_mem_counter[3007] = 4'b0000;
    GSharePlugin_logic_mem_counter[3008] = 4'b0000;
    GSharePlugin_logic_mem_counter[3009] = 4'b0000;
    GSharePlugin_logic_mem_counter[3010] = 4'b0000;
    GSharePlugin_logic_mem_counter[3011] = 4'b0000;
    GSharePlugin_logic_mem_counter[3012] = 4'b0000;
    GSharePlugin_logic_mem_counter[3013] = 4'b0000;
    GSharePlugin_logic_mem_counter[3014] = 4'b0000;
    GSharePlugin_logic_mem_counter[3015] = 4'b0000;
    GSharePlugin_logic_mem_counter[3016] = 4'b0000;
    GSharePlugin_logic_mem_counter[3017] = 4'b0000;
    GSharePlugin_logic_mem_counter[3018] = 4'b0000;
    GSharePlugin_logic_mem_counter[3019] = 4'b0000;
    GSharePlugin_logic_mem_counter[3020] = 4'b0000;
    GSharePlugin_logic_mem_counter[3021] = 4'b0000;
    GSharePlugin_logic_mem_counter[3022] = 4'b0000;
    GSharePlugin_logic_mem_counter[3023] = 4'b0000;
    GSharePlugin_logic_mem_counter[3024] = 4'b0000;
    GSharePlugin_logic_mem_counter[3025] = 4'b0000;
    GSharePlugin_logic_mem_counter[3026] = 4'b0000;
    GSharePlugin_logic_mem_counter[3027] = 4'b0000;
    GSharePlugin_logic_mem_counter[3028] = 4'b0000;
    GSharePlugin_logic_mem_counter[3029] = 4'b0000;
    GSharePlugin_logic_mem_counter[3030] = 4'b0000;
    GSharePlugin_logic_mem_counter[3031] = 4'b0000;
    GSharePlugin_logic_mem_counter[3032] = 4'b0000;
    GSharePlugin_logic_mem_counter[3033] = 4'b0000;
    GSharePlugin_logic_mem_counter[3034] = 4'b0000;
    GSharePlugin_logic_mem_counter[3035] = 4'b0000;
    GSharePlugin_logic_mem_counter[3036] = 4'b0000;
    GSharePlugin_logic_mem_counter[3037] = 4'b0000;
    GSharePlugin_logic_mem_counter[3038] = 4'b0000;
    GSharePlugin_logic_mem_counter[3039] = 4'b0000;
    GSharePlugin_logic_mem_counter[3040] = 4'b0000;
    GSharePlugin_logic_mem_counter[3041] = 4'b0000;
    GSharePlugin_logic_mem_counter[3042] = 4'b0000;
    GSharePlugin_logic_mem_counter[3043] = 4'b0000;
    GSharePlugin_logic_mem_counter[3044] = 4'b0000;
    GSharePlugin_logic_mem_counter[3045] = 4'b0000;
    GSharePlugin_logic_mem_counter[3046] = 4'b0000;
    GSharePlugin_logic_mem_counter[3047] = 4'b0000;
    GSharePlugin_logic_mem_counter[3048] = 4'b0000;
    GSharePlugin_logic_mem_counter[3049] = 4'b0000;
    GSharePlugin_logic_mem_counter[3050] = 4'b0000;
    GSharePlugin_logic_mem_counter[3051] = 4'b0000;
    GSharePlugin_logic_mem_counter[3052] = 4'b0000;
    GSharePlugin_logic_mem_counter[3053] = 4'b0000;
    GSharePlugin_logic_mem_counter[3054] = 4'b0000;
    GSharePlugin_logic_mem_counter[3055] = 4'b0000;
    GSharePlugin_logic_mem_counter[3056] = 4'b0000;
    GSharePlugin_logic_mem_counter[3057] = 4'b0000;
    GSharePlugin_logic_mem_counter[3058] = 4'b0000;
    GSharePlugin_logic_mem_counter[3059] = 4'b0000;
    GSharePlugin_logic_mem_counter[3060] = 4'b0000;
    GSharePlugin_logic_mem_counter[3061] = 4'b0000;
    GSharePlugin_logic_mem_counter[3062] = 4'b0000;
    GSharePlugin_logic_mem_counter[3063] = 4'b0000;
    GSharePlugin_logic_mem_counter[3064] = 4'b0000;
    GSharePlugin_logic_mem_counter[3065] = 4'b0000;
    GSharePlugin_logic_mem_counter[3066] = 4'b0000;
    GSharePlugin_logic_mem_counter[3067] = 4'b0000;
    GSharePlugin_logic_mem_counter[3068] = 4'b0000;
    GSharePlugin_logic_mem_counter[3069] = 4'b0000;
    GSharePlugin_logic_mem_counter[3070] = 4'b0000;
    GSharePlugin_logic_mem_counter[3071] = 4'b0000;
    GSharePlugin_logic_mem_counter[3072] = 4'b0000;
    GSharePlugin_logic_mem_counter[3073] = 4'b0000;
    GSharePlugin_logic_mem_counter[3074] = 4'b0000;
    GSharePlugin_logic_mem_counter[3075] = 4'b0000;
    GSharePlugin_logic_mem_counter[3076] = 4'b0000;
    GSharePlugin_logic_mem_counter[3077] = 4'b0000;
    GSharePlugin_logic_mem_counter[3078] = 4'b0000;
    GSharePlugin_logic_mem_counter[3079] = 4'b0000;
    GSharePlugin_logic_mem_counter[3080] = 4'b0000;
    GSharePlugin_logic_mem_counter[3081] = 4'b0000;
    GSharePlugin_logic_mem_counter[3082] = 4'b0000;
    GSharePlugin_logic_mem_counter[3083] = 4'b0000;
    GSharePlugin_logic_mem_counter[3084] = 4'b0000;
    GSharePlugin_logic_mem_counter[3085] = 4'b0000;
    GSharePlugin_logic_mem_counter[3086] = 4'b0000;
    GSharePlugin_logic_mem_counter[3087] = 4'b0000;
    GSharePlugin_logic_mem_counter[3088] = 4'b0000;
    GSharePlugin_logic_mem_counter[3089] = 4'b0000;
    GSharePlugin_logic_mem_counter[3090] = 4'b0000;
    GSharePlugin_logic_mem_counter[3091] = 4'b0000;
    GSharePlugin_logic_mem_counter[3092] = 4'b0000;
    GSharePlugin_logic_mem_counter[3093] = 4'b0000;
    GSharePlugin_logic_mem_counter[3094] = 4'b0000;
    GSharePlugin_logic_mem_counter[3095] = 4'b0000;
    GSharePlugin_logic_mem_counter[3096] = 4'b0000;
    GSharePlugin_logic_mem_counter[3097] = 4'b0000;
    GSharePlugin_logic_mem_counter[3098] = 4'b0000;
    GSharePlugin_logic_mem_counter[3099] = 4'b0000;
    GSharePlugin_logic_mem_counter[3100] = 4'b0000;
    GSharePlugin_logic_mem_counter[3101] = 4'b0000;
    GSharePlugin_logic_mem_counter[3102] = 4'b0000;
    GSharePlugin_logic_mem_counter[3103] = 4'b0000;
    GSharePlugin_logic_mem_counter[3104] = 4'b0000;
    GSharePlugin_logic_mem_counter[3105] = 4'b0000;
    GSharePlugin_logic_mem_counter[3106] = 4'b0000;
    GSharePlugin_logic_mem_counter[3107] = 4'b0000;
    GSharePlugin_logic_mem_counter[3108] = 4'b0000;
    GSharePlugin_logic_mem_counter[3109] = 4'b0000;
    GSharePlugin_logic_mem_counter[3110] = 4'b0000;
    GSharePlugin_logic_mem_counter[3111] = 4'b0000;
    GSharePlugin_logic_mem_counter[3112] = 4'b0000;
    GSharePlugin_logic_mem_counter[3113] = 4'b0000;
    GSharePlugin_logic_mem_counter[3114] = 4'b0000;
    GSharePlugin_logic_mem_counter[3115] = 4'b0000;
    GSharePlugin_logic_mem_counter[3116] = 4'b0000;
    GSharePlugin_logic_mem_counter[3117] = 4'b0000;
    GSharePlugin_logic_mem_counter[3118] = 4'b0000;
    GSharePlugin_logic_mem_counter[3119] = 4'b0000;
    GSharePlugin_logic_mem_counter[3120] = 4'b0000;
    GSharePlugin_logic_mem_counter[3121] = 4'b0000;
    GSharePlugin_logic_mem_counter[3122] = 4'b0000;
    GSharePlugin_logic_mem_counter[3123] = 4'b0000;
    GSharePlugin_logic_mem_counter[3124] = 4'b0000;
    GSharePlugin_logic_mem_counter[3125] = 4'b0000;
    GSharePlugin_logic_mem_counter[3126] = 4'b0000;
    GSharePlugin_logic_mem_counter[3127] = 4'b0000;
    GSharePlugin_logic_mem_counter[3128] = 4'b0000;
    GSharePlugin_logic_mem_counter[3129] = 4'b0000;
    GSharePlugin_logic_mem_counter[3130] = 4'b0000;
    GSharePlugin_logic_mem_counter[3131] = 4'b0000;
    GSharePlugin_logic_mem_counter[3132] = 4'b0000;
    GSharePlugin_logic_mem_counter[3133] = 4'b0000;
    GSharePlugin_logic_mem_counter[3134] = 4'b0000;
    GSharePlugin_logic_mem_counter[3135] = 4'b0000;
    GSharePlugin_logic_mem_counter[3136] = 4'b0000;
    GSharePlugin_logic_mem_counter[3137] = 4'b0000;
    GSharePlugin_logic_mem_counter[3138] = 4'b0000;
    GSharePlugin_logic_mem_counter[3139] = 4'b0000;
    GSharePlugin_logic_mem_counter[3140] = 4'b0000;
    GSharePlugin_logic_mem_counter[3141] = 4'b0000;
    GSharePlugin_logic_mem_counter[3142] = 4'b0000;
    GSharePlugin_logic_mem_counter[3143] = 4'b0000;
    GSharePlugin_logic_mem_counter[3144] = 4'b0000;
    GSharePlugin_logic_mem_counter[3145] = 4'b0000;
    GSharePlugin_logic_mem_counter[3146] = 4'b0000;
    GSharePlugin_logic_mem_counter[3147] = 4'b0000;
    GSharePlugin_logic_mem_counter[3148] = 4'b0000;
    GSharePlugin_logic_mem_counter[3149] = 4'b0000;
    GSharePlugin_logic_mem_counter[3150] = 4'b0000;
    GSharePlugin_logic_mem_counter[3151] = 4'b0000;
    GSharePlugin_logic_mem_counter[3152] = 4'b0000;
    GSharePlugin_logic_mem_counter[3153] = 4'b0000;
    GSharePlugin_logic_mem_counter[3154] = 4'b0000;
    GSharePlugin_logic_mem_counter[3155] = 4'b0000;
    GSharePlugin_logic_mem_counter[3156] = 4'b0000;
    GSharePlugin_logic_mem_counter[3157] = 4'b0000;
    GSharePlugin_logic_mem_counter[3158] = 4'b0000;
    GSharePlugin_logic_mem_counter[3159] = 4'b0000;
    GSharePlugin_logic_mem_counter[3160] = 4'b0000;
    GSharePlugin_logic_mem_counter[3161] = 4'b0000;
    GSharePlugin_logic_mem_counter[3162] = 4'b0000;
    GSharePlugin_logic_mem_counter[3163] = 4'b0000;
    GSharePlugin_logic_mem_counter[3164] = 4'b0000;
    GSharePlugin_logic_mem_counter[3165] = 4'b0000;
    GSharePlugin_logic_mem_counter[3166] = 4'b0000;
    GSharePlugin_logic_mem_counter[3167] = 4'b0000;
    GSharePlugin_logic_mem_counter[3168] = 4'b0000;
    GSharePlugin_logic_mem_counter[3169] = 4'b0000;
    GSharePlugin_logic_mem_counter[3170] = 4'b0000;
    GSharePlugin_logic_mem_counter[3171] = 4'b0000;
    GSharePlugin_logic_mem_counter[3172] = 4'b0000;
    GSharePlugin_logic_mem_counter[3173] = 4'b0000;
    GSharePlugin_logic_mem_counter[3174] = 4'b0000;
    GSharePlugin_logic_mem_counter[3175] = 4'b0000;
    GSharePlugin_logic_mem_counter[3176] = 4'b0000;
    GSharePlugin_logic_mem_counter[3177] = 4'b0000;
    GSharePlugin_logic_mem_counter[3178] = 4'b0000;
    GSharePlugin_logic_mem_counter[3179] = 4'b0000;
    GSharePlugin_logic_mem_counter[3180] = 4'b0000;
    GSharePlugin_logic_mem_counter[3181] = 4'b0000;
    GSharePlugin_logic_mem_counter[3182] = 4'b0000;
    GSharePlugin_logic_mem_counter[3183] = 4'b0000;
    GSharePlugin_logic_mem_counter[3184] = 4'b0000;
    GSharePlugin_logic_mem_counter[3185] = 4'b0000;
    GSharePlugin_logic_mem_counter[3186] = 4'b0000;
    GSharePlugin_logic_mem_counter[3187] = 4'b0000;
    GSharePlugin_logic_mem_counter[3188] = 4'b0000;
    GSharePlugin_logic_mem_counter[3189] = 4'b0000;
    GSharePlugin_logic_mem_counter[3190] = 4'b0000;
    GSharePlugin_logic_mem_counter[3191] = 4'b0000;
    GSharePlugin_logic_mem_counter[3192] = 4'b0000;
    GSharePlugin_logic_mem_counter[3193] = 4'b0000;
    GSharePlugin_logic_mem_counter[3194] = 4'b0000;
    GSharePlugin_logic_mem_counter[3195] = 4'b0000;
    GSharePlugin_logic_mem_counter[3196] = 4'b0000;
    GSharePlugin_logic_mem_counter[3197] = 4'b0000;
    GSharePlugin_logic_mem_counter[3198] = 4'b0000;
    GSharePlugin_logic_mem_counter[3199] = 4'b0000;
    GSharePlugin_logic_mem_counter[3200] = 4'b0000;
    GSharePlugin_logic_mem_counter[3201] = 4'b0000;
    GSharePlugin_logic_mem_counter[3202] = 4'b0000;
    GSharePlugin_logic_mem_counter[3203] = 4'b0000;
    GSharePlugin_logic_mem_counter[3204] = 4'b0000;
    GSharePlugin_logic_mem_counter[3205] = 4'b0000;
    GSharePlugin_logic_mem_counter[3206] = 4'b0000;
    GSharePlugin_logic_mem_counter[3207] = 4'b0000;
    GSharePlugin_logic_mem_counter[3208] = 4'b0000;
    GSharePlugin_logic_mem_counter[3209] = 4'b0000;
    GSharePlugin_logic_mem_counter[3210] = 4'b0000;
    GSharePlugin_logic_mem_counter[3211] = 4'b0000;
    GSharePlugin_logic_mem_counter[3212] = 4'b0000;
    GSharePlugin_logic_mem_counter[3213] = 4'b0000;
    GSharePlugin_logic_mem_counter[3214] = 4'b0000;
    GSharePlugin_logic_mem_counter[3215] = 4'b0000;
    GSharePlugin_logic_mem_counter[3216] = 4'b0000;
    GSharePlugin_logic_mem_counter[3217] = 4'b0000;
    GSharePlugin_logic_mem_counter[3218] = 4'b0000;
    GSharePlugin_logic_mem_counter[3219] = 4'b0000;
    GSharePlugin_logic_mem_counter[3220] = 4'b0000;
    GSharePlugin_logic_mem_counter[3221] = 4'b0000;
    GSharePlugin_logic_mem_counter[3222] = 4'b0000;
    GSharePlugin_logic_mem_counter[3223] = 4'b0000;
    GSharePlugin_logic_mem_counter[3224] = 4'b0000;
    GSharePlugin_logic_mem_counter[3225] = 4'b0000;
    GSharePlugin_logic_mem_counter[3226] = 4'b0000;
    GSharePlugin_logic_mem_counter[3227] = 4'b0000;
    GSharePlugin_logic_mem_counter[3228] = 4'b0000;
    GSharePlugin_logic_mem_counter[3229] = 4'b0000;
    GSharePlugin_logic_mem_counter[3230] = 4'b0000;
    GSharePlugin_logic_mem_counter[3231] = 4'b0000;
    GSharePlugin_logic_mem_counter[3232] = 4'b0000;
    GSharePlugin_logic_mem_counter[3233] = 4'b0000;
    GSharePlugin_logic_mem_counter[3234] = 4'b0000;
    GSharePlugin_logic_mem_counter[3235] = 4'b0000;
    GSharePlugin_logic_mem_counter[3236] = 4'b0000;
    GSharePlugin_logic_mem_counter[3237] = 4'b0000;
    GSharePlugin_logic_mem_counter[3238] = 4'b0000;
    GSharePlugin_logic_mem_counter[3239] = 4'b0000;
    GSharePlugin_logic_mem_counter[3240] = 4'b0000;
    GSharePlugin_logic_mem_counter[3241] = 4'b0000;
    GSharePlugin_logic_mem_counter[3242] = 4'b0000;
    GSharePlugin_logic_mem_counter[3243] = 4'b0000;
    GSharePlugin_logic_mem_counter[3244] = 4'b0000;
    GSharePlugin_logic_mem_counter[3245] = 4'b0000;
    GSharePlugin_logic_mem_counter[3246] = 4'b0000;
    GSharePlugin_logic_mem_counter[3247] = 4'b0000;
    GSharePlugin_logic_mem_counter[3248] = 4'b0000;
    GSharePlugin_logic_mem_counter[3249] = 4'b0000;
    GSharePlugin_logic_mem_counter[3250] = 4'b0000;
    GSharePlugin_logic_mem_counter[3251] = 4'b0000;
    GSharePlugin_logic_mem_counter[3252] = 4'b0000;
    GSharePlugin_logic_mem_counter[3253] = 4'b0000;
    GSharePlugin_logic_mem_counter[3254] = 4'b0000;
    GSharePlugin_logic_mem_counter[3255] = 4'b0000;
    GSharePlugin_logic_mem_counter[3256] = 4'b0000;
    GSharePlugin_logic_mem_counter[3257] = 4'b0000;
    GSharePlugin_logic_mem_counter[3258] = 4'b0000;
    GSharePlugin_logic_mem_counter[3259] = 4'b0000;
    GSharePlugin_logic_mem_counter[3260] = 4'b0000;
    GSharePlugin_logic_mem_counter[3261] = 4'b0000;
    GSharePlugin_logic_mem_counter[3262] = 4'b0000;
    GSharePlugin_logic_mem_counter[3263] = 4'b0000;
    GSharePlugin_logic_mem_counter[3264] = 4'b0000;
    GSharePlugin_logic_mem_counter[3265] = 4'b0000;
    GSharePlugin_logic_mem_counter[3266] = 4'b0000;
    GSharePlugin_logic_mem_counter[3267] = 4'b0000;
    GSharePlugin_logic_mem_counter[3268] = 4'b0000;
    GSharePlugin_logic_mem_counter[3269] = 4'b0000;
    GSharePlugin_logic_mem_counter[3270] = 4'b0000;
    GSharePlugin_logic_mem_counter[3271] = 4'b0000;
    GSharePlugin_logic_mem_counter[3272] = 4'b0000;
    GSharePlugin_logic_mem_counter[3273] = 4'b0000;
    GSharePlugin_logic_mem_counter[3274] = 4'b0000;
    GSharePlugin_logic_mem_counter[3275] = 4'b0000;
    GSharePlugin_logic_mem_counter[3276] = 4'b0000;
    GSharePlugin_logic_mem_counter[3277] = 4'b0000;
    GSharePlugin_logic_mem_counter[3278] = 4'b0000;
    GSharePlugin_logic_mem_counter[3279] = 4'b0000;
    GSharePlugin_logic_mem_counter[3280] = 4'b0000;
    GSharePlugin_logic_mem_counter[3281] = 4'b0000;
    GSharePlugin_logic_mem_counter[3282] = 4'b0000;
    GSharePlugin_logic_mem_counter[3283] = 4'b0000;
    GSharePlugin_logic_mem_counter[3284] = 4'b0000;
    GSharePlugin_logic_mem_counter[3285] = 4'b0000;
    GSharePlugin_logic_mem_counter[3286] = 4'b0000;
    GSharePlugin_logic_mem_counter[3287] = 4'b0000;
    GSharePlugin_logic_mem_counter[3288] = 4'b0000;
    GSharePlugin_logic_mem_counter[3289] = 4'b0000;
    GSharePlugin_logic_mem_counter[3290] = 4'b0000;
    GSharePlugin_logic_mem_counter[3291] = 4'b0000;
    GSharePlugin_logic_mem_counter[3292] = 4'b0000;
    GSharePlugin_logic_mem_counter[3293] = 4'b0000;
    GSharePlugin_logic_mem_counter[3294] = 4'b0000;
    GSharePlugin_logic_mem_counter[3295] = 4'b0000;
    GSharePlugin_logic_mem_counter[3296] = 4'b0000;
    GSharePlugin_logic_mem_counter[3297] = 4'b0000;
    GSharePlugin_logic_mem_counter[3298] = 4'b0000;
    GSharePlugin_logic_mem_counter[3299] = 4'b0000;
    GSharePlugin_logic_mem_counter[3300] = 4'b0000;
    GSharePlugin_logic_mem_counter[3301] = 4'b0000;
    GSharePlugin_logic_mem_counter[3302] = 4'b0000;
    GSharePlugin_logic_mem_counter[3303] = 4'b0000;
    GSharePlugin_logic_mem_counter[3304] = 4'b0000;
    GSharePlugin_logic_mem_counter[3305] = 4'b0000;
    GSharePlugin_logic_mem_counter[3306] = 4'b0000;
    GSharePlugin_logic_mem_counter[3307] = 4'b0000;
    GSharePlugin_logic_mem_counter[3308] = 4'b0000;
    GSharePlugin_logic_mem_counter[3309] = 4'b0000;
    GSharePlugin_logic_mem_counter[3310] = 4'b0000;
    GSharePlugin_logic_mem_counter[3311] = 4'b0000;
    GSharePlugin_logic_mem_counter[3312] = 4'b0000;
    GSharePlugin_logic_mem_counter[3313] = 4'b0000;
    GSharePlugin_logic_mem_counter[3314] = 4'b0000;
    GSharePlugin_logic_mem_counter[3315] = 4'b0000;
    GSharePlugin_logic_mem_counter[3316] = 4'b0000;
    GSharePlugin_logic_mem_counter[3317] = 4'b0000;
    GSharePlugin_logic_mem_counter[3318] = 4'b0000;
    GSharePlugin_logic_mem_counter[3319] = 4'b0000;
    GSharePlugin_logic_mem_counter[3320] = 4'b0000;
    GSharePlugin_logic_mem_counter[3321] = 4'b0000;
    GSharePlugin_logic_mem_counter[3322] = 4'b0000;
    GSharePlugin_logic_mem_counter[3323] = 4'b0000;
    GSharePlugin_logic_mem_counter[3324] = 4'b0000;
    GSharePlugin_logic_mem_counter[3325] = 4'b0000;
    GSharePlugin_logic_mem_counter[3326] = 4'b0000;
    GSharePlugin_logic_mem_counter[3327] = 4'b0000;
    GSharePlugin_logic_mem_counter[3328] = 4'b0000;
    GSharePlugin_logic_mem_counter[3329] = 4'b0000;
    GSharePlugin_logic_mem_counter[3330] = 4'b0000;
    GSharePlugin_logic_mem_counter[3331] = 4'b0000;
    GSharePlugin_logic_mem_counter[3332] = 4'b0000;
    GSharePlugin_logic_mem_counter[3333] = 4'b0000;
    GSharePlugin_logic_mem_counter[3334] = 4'b0000;
    GSharePlugin_logic_mem_counter[3335] = 4'b0000;
    GSharePlugin_logic_mem_counter[3336] = 4'b0000;
    GSharePlugin_logic_mem_counter[3337] = 4'b0000;
    GSharePlugin_logic_mem_counter[3338] = 4'b0000;
    GSharePlugin_logic_mem_counter[3339] = 4'b0000;
    GSharePlugin_logic_mem_counter[3340] = 4'b0000;
    GSharePlugin_logic_mem_counter[3341] = 4'b0000;
    GSharePlugin_logic_mem_counter[3342] = 4'b0000;
    GSharePlugin_logic_mem_counter[3343] = 4'b0000;
    GSharePlugin_logic_mem_counter[3344] = 4'b0000;
    GSharePlugin_logic_mem_counter[3345] = 4'b0000;
    GSharePlugin_logic_mem_counter[3346] = 4'b0000;
    GSharePlugin_logic_mem_counter[3347] = 4'b0000;
    GSharePlugin_logic_mem_counter[3348] = 4'b0000;
    GSharePlugin_logic_mem_counter[3349] = 4'b0000;
    GSharePlugin_logic_mem_counter[3350] = 4'b0000;
    GSharePlugin_logic_mem_counter[3351] = 4'b0000;
    GSharePlugin_logic_mem_counter[3352] = 4'b0000;
    GSharePlugin_logic_mem_counter[3353] = 4'b0000;
    GSharePlugin_logic_mem_counter[3354] = 4'b0000;
    GSharePlugin_logic_mem_counter[3355] = 4'b0000;
    GSharePlugin_logic_mem_counter[3356] = 4'b0000;
    GSharePlugin_logic_mem_counter[3357] = 4'b0000;
    GSharePlugin_logic_mem_counter[3358] = 4'b0000;
    GSharePlugin_logic_mem_counter[3359] = 4'b0000;
    GSharePlugin_logic_mem_counter[3360] = 4'b0000;
    GSharePlugin_logic_mem_counter[3361] = 4'b0000;
    GSharePlugin_logic_mem_counter[3362] = 4'b0000;
    GSharePlugin_logic_mem_counter[3363] = 4'b0000;
    GSharePlugin_logic_mem_counter[3364] = 4'b0000;
    GSharePlugin_logic_mem_counter[3365] = 4'b0000;
    GSharePlugin_logic_mem_counter[3366] = 4'b0000;
    GSharePlugin_logic_mem_counter[3367] = 4'b0000;
    GSharePlugin_logic_mem_counter[3368] = 4'b0000;
    GSharePlugin_logic_mem_counter[3369] = 4'b0000;
    GSharePlugin_logic_mem_counter[3370] = 4'b0000;
    GSharePlugin_logic_mem_counter[3371] = 4'b0000;
    GSharePlugin_logic_mem_counter[3372] = 4'b0000;
    GSharePlugin_logic_mem_counter[3373] = 4'b0000;
    GSharePlugin_logic_mem_counter[3374] = 4'b0000;
    GSharePlugin_logic_mem_counter[3375] = 4'b0000;
    GSharePlugin_logic_mem_counter[3376] = 4'b0000;
    GSharePlugin_logic_mem_counter[3377] = 4'b0000;
    GSharePlugin_logic_mem_counter[3378] = 4'b0000;
    GSharePlugin_logic_mem_counter[3379] = 4'b0000;
    GSharePlugin_logic_mem_counter[3380] = 4'b0000;
    GSharePlugin_logic_mem_counter[3381] = 4'b0000;
    GSharePlugin_logic_mem_counter[3382] = 4'b0000;
    GSharePlugin_logic_mem_counter[3383] = 4'b0000;
    GSharePlugin_logic_mem_counter[3384] = 4'b0000;
    GSharePlugin_logic_mem_counter[3385] = 4'b0000;
    GSharePlugin_logic_mem_counter[3386] = 4'b0000;
    GSharePlugin_logic_mem_counter[3387] = 4'b0000;
    GSharePlugin_logic_mem_counter[3388] = 4'b0000;
    GSharePlugin_logic_mem_counter[3389] = 4'b0000;
    GSharePlugin_logic_mem_counter[3390] = 4'b0000;
    GSharePlugin_logic_mem_counter[3391] = 4'b0000;
    GSharePlugin_logic_mem_counter[3392] = 4'b0000;
    GSharePlugin_logic_mem_counter[3393] = 4'b0000;
    GSharePlugin_logic_mem_counter[3394] = 4'b0000;
    GSharePlugin_logic_mem_counter[3395] = 4'b0000;
    GSharePlugin_logic_mem_counter[3396] = 4'b0000;
    GSharePlugin_logic_mem_counter[3397] = 4'b0000;
    GSharePlugin_logic_mem_counter[3398] = 4'b0000;
    GSharePlugin_logic_mem_counter[3399] = 4'b0000;
    GSharePlugin_logic_mem_counter[3400] = 4'b0000;
    GSharePlugin_logic_mem_counter[3401] = 4'b0000;
    GSharePlugin_logic_mem_counter[3402] = 4'b0000;
    GSharePlugin_logic_mem_counter[3403] = 4'b0000;
    GSharePlugin_logic_mem_counter[3404] = 4'b0000;
    GSharePlugin_logic_mem_counter[3405] = 4'b0000;
    GSharePlugin_logic_mem_counter[3406] = 4'b0000;
    GSharePlugin_logic_mem_counter[3407] = 4'b0000;
    GSharePlugin_logic_mem_counter[3408] = 4'b0000;
    GSharePlugin_logic_mem_counter[3409] = 4'b0000;
    GSharePlugin_logic_mem_counter[3410] = 4'b0000;
    GSharePlugin_logic_mem_counter[3411] = 4'b0000;
    GSharePlugin_logic_mem_counter[3412] = 4'b0000;
    GSharePlugin_logic_mem_counter[3413] = 4'b0000;
    GSharePlugin_logic_mem_counter[3414] = 4'b0000;
    GSharePlugin_logic_mem_counter[3415] = 4'b0000;
    GSharePlugin_logic_mem_counter[3416] = 4'b0000;
    GSharePlugin_logic_mem_counter[3417] = 4'b0000;
    GSharePlugin_logic_mem_counter[3418] = 4'b0000;
    GSharePlugin_logic_mem_counter[3419] = 4'b0000;
    GSharePlugin_logic_mem_counter[3420] = 4'b0000;
    GSharePlugin_logic_mem_counter[3421] = 4'b0000;
    GSharePlugin_logic_mem_counter[3422] = 4'b0000;
    GSharePlugin_logic_mem_counter[3423] = 4'b0000;
    GSharePlugin_logic_mem_counter[3424] = 4'b0000;
    GSharePlugin_logic_mem_counter[3425] = 4'b0000;
    GSharePlugin_logic_mem_counter[3426] = 4'b0000;
    GSharePlugin_logic_mem_counter[3427] = 4'b0000;
    GSharePlugin_logic_mem_counter[3428] = 4'b0000;
    GSharePlugin_logic_mem_counter[3429] = 4'b0000;
    GSharePlugin_logic_mem_counter[3430] = 4'b0000;
    GSharePlugin_logic_mem_counter[3431] = 4'b0000;
    GSharePlugin_logic_mem_counter[3432] = 4'b0000;
    GSharePlugin_logic_mem_counter[3433] = 4'b0000;
    GSharePlugin_logic_mem_counter[3434] = 4'b0000;
    GSharePlugin_logic_mem_counter[3435] = 4'b0000;
    GSharePlugin_logic_mem_counter[3436] = 4'b0000;
    GSharePlugin_logic_mem_counter[3437] = 4'b0000;
    GSharePlugin_logic_mem_counter[3438] = 4'b0000;
    GSharePlugin_logic_mem_counter[3439] = 4'b0000;
    GSharePlugin_logic_mem_counter[3440] = 4'b0000;
    GSharePlugin_logic_mem_counter[3441] = 4'b0000;
    GSharePlugin_logic_mem_counter[3442] = 4'b0000;
    GSharePlugin_logic_mem_counter[3443] = 4'b0000;
    GSharePlugin_logic_mem_counter[3444] = 4'b0000;
    GSharePlugin_logic_mem_counter[3445] = 4'b0000;
    GSharePlugin_logic_mem_counter[3446] = 4'b0000;
    GSharePlugin_logic_mem_counter[3447] = 4'b0000;
    GSharePlugin_logic_mem_counter[3448] = 4'b0000;
    GSharePlugin_logic_mem_counter[3449] = 4'b0000;
    GSharePlugin_logic_mem_counter[3450] = 4'b0000;
    GSharePlugin_logic_mem_counter[3451] = 4'b0000;
    GSharePlugin_logic_mem_counter[3452] = 4'b0000;
    GSharePlugin_logic_mem_counter[3453] = 4'b0000;
    GSharePlugin_logic_mem_counter[3454] = 4'b0000;
    GSharePlugin_logic_mem_counter[3455] = 4'b0000;
    GSharePlugin_logic_mem_counter[3456] = 4'b0000;
    GSharePlugin_logic_mem_counter[3457] = 4'b0000;
    GSharePlugin_logic_mem_counter[3458] = 4'b0000;
    GSharePlugin_logic_mem_counter[3459] = 4'b0000;
    GSharePlugin_logic_mem_counter[3460] = 4'b0000;
    GSharePlugin_logic_mem_counter[3461] = 4'b0000;
    GSharePlugin_logic_mem_counter[3462] = 4'b0000;
    GSharePlugin_logic_mem_counter[3463] = 4'b0000;
    GSharePlugin_logic_mem_counter[3464] = 4'b0000;
    GSharePlugin_logic_mem_counter[3465] = 4'b0000;
    GSharePlugin_logic_mem_counter[3466] = 4'b0000;
    GSharePlugin_logic_mem_counter[3467] = 4'b0000;
    GSharePlugin_logic_mem_counter[3468] = 4'b0000;
    GSharePlugin_logic_mem_counter[3469] = 4'b0000;
    GSharePlugin_logic_mem_counter[3470] = 4'b0000;
    GSharePlugin_logic_mem_counter[3471] = 4'b0000;
    GSharePlugin_logic_mem_counter[3472] = 4'b0000;
    GSharePlugin_logic_mem_counter[3473] = 4'b0000;
    GSharePlugin_logic_mem_counter[3474] = 4'b0000;
    GSharePlugin_logic_mem_counter[3475] = 4'b0000;
    GSharePlugin_logic_mem_counter[3476] = 4'b0000;
    GSharePlugin_logic_mem_counter[3477] = 4'b0000;
    GSharePlugin_logic_mem_counter[3478] = 4'b0000;
    GSharePlugin_logic_mem_counter[3479] = 4'b0000;
    GSharePlugin_logic_mem_counter[3480] = 4'b0000;
    GSharePlugin_logic_mem_counter[3481] = 4'b0000;
    GSharePlugin_logic_mem_counter[3482] = 4'b0000;
    GSharePlugin_logic_mem_counter[3483] = 4'b0000;
    GSharePlugin_logic_mem_counter[3484] = 4'b0000;
    GSharePlugin_logic_mem_counter[3485] = 4'b0000;
    GSharePlugin_logic_mem_counter[3486] = 4'b0000;
    GSharePlugin_logic_mem_counter[3487] = 4'b0000;
    GSharePlugin_logic_mem_counter[3488] = 4'b0000;
    GSharePlugin_logic_mem_counter[3489] = 4'b0000;
    GSharePlugin_logic_mem_counter[3490] = 4'b0000;
    GSharePlugin_logic_mem_counter[3491] = 4'b0000;
    GSharePlugin_logic_mem_counter[3492] = 4'b0000;
    GSharePlugin_logic_mem_counter[3493] = 4'b0000;
    GSharePlugin_logic_mem_counter[3494] = 4'b0000;
    GSharePlugin_logic_mem_counter[3495] = 4'b0000;
    GSharePlugin_logic_mem_counter[3496] = 4'b0000;
    GSharePlugin_logic_mem_counter[3497] = 4'b0000;
    GSharePlugin_logic_mem_counter[3498] = 4'b0000;
    GSharePlugin_logic_mem_counter[3499] = 4'b0000;
    GSharePlugin_logic_mem_counter[3500] = 4'b0000;
    GSharePlugin_logic_mem_counter[3501] = 4'b0000;
    GSharePlugin_logic_mem_counter[3502] = 4'b0000;
    GSharePlugin_logic_mem_counter[3503] = 4'b0000;
    GSharePlugin_logic_mem_counter[3504] = 4'b0000;
    GSharePlugin_logic_mem_counter[3505] = 4'b0000;
    GSharePlugin_logic_mem_counter[3506] = 4'b0000;
    GSharePlugin_logic_mem_counter[3507] = 4'b0000;
    GSharePlugin_logic_mem_counter[3508] = 4'b0000;
    GSharePlugin_logic_mem_counter[3509] = 4'b0000;
    GSharePlugin_logic_mem_counter[3510] = 4'b0000;
    GSharePlugin_logic_mem_counter[3511] = 4'b0000;
    GSharePlugin_logic_mem_counter[3512] = 4'b0000;
    GSharePlugin_logic_mem_counter[3513] = 4'b0000;
    GSharePlugin_logic_mem_counter[3514] = 4'b0000;
    GSharePlugin_logic_mem_counter[3515] = 4'b0000;
    GSharePlugin_logic_mem_counter[3516] = 4'b0000;
    GSharePlugin_logic_mem_counter[3517] = 4'b0000;
    GSharePlugin_logic_mem_counter[3518] = 4'b0000;
    GSharePlugin_logic_mem_counter[3519] = 4'b0000;
    GSharePlugin_logic_mem_counter[3520] = 4'b0000;
    GSharePlugin_logic_mem_counter[3521] = 4'b0000;
    GSharePlugin_logic_mem_counter[3522] = 4'b0000;
    GSharePlugin_logic_mem_counter[3523] = 4'b0000;
    GSharePlugin_logic_mem_counter[3524] = 4'b0000;
    GSharePlugin_logic_mem_counter[3525] = 4'b0000;
    GSharePlugin_logic_mem_counter[3526] = 4'b0000;
    GSharePlugin_logic_mem_counter[3527] = 4'b0000;
    GSharePlugin_logic_mem_counter[3528] = 4'b0000;
    GSharePlugin_logic_mem_counter[3529] = 4'b0000;
    GSharePlugin_logic_mem_counter[3530] = 4'b0000;
    GSharePlugin_logic_mem_counter[3531] = 4'b0000;
    GSharePlugin_logic_mem_counter[3532] = 4'b0000;
    GSharePlugin_logic_mem_counter[3533] = 4'b0000;
    GSharePlugin_logic_mem_counter[3534] = 4'b0000;
    GSharePlugin_logic_mem_counter[3535] = 4'b0000;
    GSharePlugin_logic_mem_counter[3536] = 4'b0000;
    GSharePlugin_logic_mem_counter[3537] = 4'b0000;
    GSharePlugin_logic_mem_counter[3538] = 4'b0000;
    GSharePlugin_logic_mem_counter[3539] = 4'b0000;
    GSharePlugin_logic_mem_counter[3540] = 4'b0000;
    GSharePlugin_logic_mem_counter[3541] = 4'b0000;
    GSharePlugin_logic_mem_counter[3542] = 4'b0000;
    GSharePlugin_logic_mem_counter[3543] = 4'b0000;
    GSharePlugin_logic_mem_counter[3544] = 4'b0000;
    GSharePlugin_logic_mem_counter[3545] = 4'b0000;
    GSharePlugin_logic_mem_counter[3546] = 4'b0000;
    GSharePlugin_logic_mem_counter[3547] = 4'b0000;
    GSharePlugin_logic_mem_counter[3548] = 4'b0000;
    GSharePlugin_logic_mem_counter[3549] = 4'b0000;
    GSharePlugin_logic_mem_counter[3550] = 4'b0000;
    GSharePlugin_logic_mem_counter[3551] = 4'b0000;
    GSharePlugin_logic_mem_counter[3552] = 4'b0000;
    GSharePlugin_logic_mem_counter[3553] = 4'b0000;
    GSharePlugin_logic_mem_counter[3554] = 4'b0000;
    GSharePlugin_logic_mem_counter[3555] = 4'b0000;
    GSharePlugin_logic_mem_counter[3556] = 4'b0000;
    GSharePlugin_logic_mem_counter[3557] = 4'b0000;
    GSharePlugin_logic_mem_counter[3558] = 4'b0000;
    GSharePlugin_logic_mem_counter[3559] = 4'b0000;
    GSharePlugin_logic_mem_counter[3560] = 4'b0000;
    GSharePlugin_logic_mem_counter[3561] = 4'b0000;
    GSharePlugin_logic_mem_counter[3562] = 4'b0000;
    GSharePlugin_logic_mem_counter[3563] = 4'b0000;
    GSharePlugin_logic_mem_counter[3564] = 4'b0000;
    GSharePlugin_logic_mem_counter[3565] = 4'b0000;
    GSharePlugin_logic_mem_counter[3566] = 4'b0000;
    GSharePlugin_logic_mem_counter[3567] = 4'b0000;
    GSharePlugin_logic_mem_counter[3568] = 4'b0000;
    GSharePlugin_logic_mem_counter[3569] = 4'b0000;
    GSharePlugin_logic_mem_counter[3570] = 4'b0000;
    GSharePlugin_logic_mem_counter[3571] = 4'b0000;
    GSharePlugin_logic_mem_counter[3572] = 4'b0000;
    GSharePlugin_logic_mem_counter[3573] = 4'b0000;
    GSharePlugin_logic_mem_counter[3574] = 4'b0000;
    GSharePlugin_logic_mem_counter[3575] = 4'b0000;
    GSharePlugin_logic_mem_counter[3576] = 4'b0000;
    GSharePlugin_logic_mem_counter[3577] = 4'b0000;
    GSharePlugin_logic_mem_counter[3578] = 4'b0000;
    GSharePlugin_logic_mem_counter[3579] = 4'b0000;
    GSharePlugin_logic_mem_counter[3580] = 4'b0000;
    GSharePlugin_logic_mem_counter[3581] = 4'b0000;
    GSharePlugin_logic_mem_counter[3582] = 4'b0000;
    GSharePlugin_logic_mem_counter[3583] = 4'b0000;
    GSharePlugin_logic_mem_counter[3584] = 4'b0000;
    GSharePlugin_logic_mem_counter[3585] = 4'b0000;
    GSharePlugin_logic_mem_counter[3586] = 4'b0000;
    GSharePlugin_logic_mem_counter[3587] = 4'b0000;
    GSharePlugin_logic_mem_counter[3588] = 4'b0000;
    GSharePlugin_logic_mem_counter[3589] = 4'b0000;
    GSharePlugin_logic_mem_counter[3590] = 4'b0000;
    GSharePlugin_logic_mem_counter[3591] = 4'b0000;
    GSharePlugin_logic_mem_counter[3592] = 4'b0000;
    GSharePlugin_logic_mem_counter[3593] = 4'b0000;
    GSharePlugin_logic_mem_counter[3594] = 4'b0000;
    GSharePlugin_logic_mem_counter[3595] = 4'b0000;
    GSharePlugin_logic_mem_counter[3596] = 4'b0000;
    GSharePlugin_logic_mem_counter[3597] = 4'b0000;
    GSharePlugin_logic_mem_counter[3598] = 4'b0000;
    GSharePlugin_logic_mem_counter[3599] = 4'b0000;
    GSharePlugin_logic_mem_counter[3600] = 4'b0000;
    GSharePlugin_logic_mem_counter[3601] = 4'b0000;
    GSharePlugin_logic_mem_counter[3602] = 4'b0000;
    GSharePlugin_logic_mem_counter[3603] = 4'b0000;
    GSharePlugin_logic_mem_counter[3604] = 4'b0000;
    GSharePlugin_logic_mem_counter[3605] = 4'b0000;
    GSharePlugin_logic_mem_counter[3606] = 4'b0000;
    GSharePlugin_logic_mem_counter[3607] = 4'b0000;
    GSharePlugin_logic_mem_counter[3608] = 4'b0000;
    GSharePlugin_logic_mem_counter[3609] = 4'b0000;
    GSharePlugin_logic_mem_counter[3610] = 4'b0000;
    GSharePlugin_logic_mem_counter[3611] = 4'b0000;
    GSharePlugin_logic_mem_counter[3612] = 4'b0000;
    GSharePlugin_logic_mem_counter[3613] = 4'b0000;
    GSharePlugin_logic_mem_counter[3614] = 4'b0000;
    GSharePlugin_logic_mem_counter[3615] = 4'b0000;
    GSharePlugin_logic_mem_counter[3616] = 4'b0000;
    GSharePlugin_logic_mem_counter[3617] = 4'b0000;
    GSharePlugin_logic_mem_counter[3618] = 4'b0000;
    GSharePlugin_logic_mem_counter[3619] = 4'b0000;
    GSharePlugin_logic_mem_counter[3620] = 4'b0000;
    GSharePlugin_logic_mem_counter[3621] = 4'b0000;
    GSharePlugin_logic_mem_counter[3622] = 4'b0000;
    GSharePlugin_logic_mem_counter[3623] = 4'b0000;
    GSharePlugin_logic_mem_counter[3624] = 4'b0000;
    GSharePlugin_logic_mem_counter[3625] = 4'b0000;
    GSharePlugin_logic_mem_counter[3626] = 4'b0000;
    GSharePlugin_logic_mem_counter[3627] = 4'b0000;
    GSharePlugin_logic_mem_counter[3628] = 4'b0000;
    GSharePlugin_logic_mem_counter[3629] = 4'b0000;
    GSharePlugin_logic_mem_counter[3630] = 4'b0000;
    GSharePlugin_logic_mem_counter[3631] = 4'b0000;
    GSharePlugin_logic_mem_counter[3632] = 4'b0000;
    GSharePlugin_logic_mem_counter[3633] = 4'b0000;
    GSharePlugin_logic_mem_counter[3634] = 4'b0000;
    GSharePlugin_logic_mem_counter[3635] = 4'b0000;
    GSharePlugin_logic_mem_counter[3636] = 4'b0000;
    GSharePlugin_logic_mem_counter[3637] = 4'b0000;
    GSharePlugin_logic_mem_counter[3638] = 4'b0000;
    GSharePlugin_logic_mem_counter[3639] = 4'b0000;
    GSharePlugin_logic_mem_counter[3640] = 4'b0000;
    GSharePlugin_logic_mem_counter[3641] = 4'b0000;
    GSharePlugin_logic_mem_counter[3642] = 4'b0000;
    GSharePlugin_logic_mem_counter[3643] = 4'b0000;
    GSharePlugin_logic_mem_counter[3644] = 4'b0000;
    GSharePlugin_logic_mem_counter[3645] = 4'b0000;
    GSharePlugin_logic_mem_counter[3646] = 4'b0000;
    GSharePlugin_logic_mem_counter[3647] = 4'b0000;
    GSharePlugin_logic_mem_counter[3648] = 4'b0000;
    GSharePlugin_logic_mem_counter[3649] = 4'b0000;
    GSharePlugin_logic_mem_counter[3650] = 4'b0000;
    GSharePlugin_logic_mem_counter[3651] = 4'b0000;
    GSharePlugin_logic_mem_counter[3652] = 4'b0000;
    GSharePlugin_logic_mem_counter[3653] = 4'b0000;
    GSharePlugin_logic_mem_counter[3654] = 4'b0000;
    GSharePlugin_logic_mem_counter[3655] = 4'b0000;
    GSharePlugin_logic_mem_counter[3656] = 4'b0000;
    GSharePlugin_logic_mem_counter[3657] = 4'b0000;
    GSharePlugin_logic_mem_counter[3658] = 4'b0000;
    GSharePlugin_logic_mem_counter[3659] = 4'b0000;
    GSharePlugin_logic_mem_counter[3660] = 4'b0000;
    GSharePlugin_logic_mem_counter[3661] = 4'b0000;
    GSharePlugin_logic_mem_counter[3662] = 4'b0000;
    GSharePlugin_logic_mem_counter[3663] = 4'b0000;
    GSharePlugin_logic_mem_counter[3664] = 4'b0000;
    GSharePlugin_logic_mem_counter[3665] = 4'b0000;
    GSharePlugin_logic_mem_counter[3666] = 4'b0000;
    GSharePlugin_logic_mem_counter[3667] = 4'b0000;
    GSharePlugin_logic_mem_counter[3668] = 4'b0000;
    GSharePlugin_logic_mem_counter[3669] = 4'b0000;
    GSharePlugin_logic_mem_counter[3670] = 4'b0000;
    GSharePlugin_logic_mem_counter[3671] = 4'b0000;
    GSharePlugin_logic_mem_counter[3672] = 4'b0000;
    GSharePlugin_logic_mem_counter[3673] = 4'b0000;
    GSharePlugin_logic_mem_counter[3674] = 4'b0000;
    GSharePlugin_logic_mem_counter[3675] = 4'b0000;
    GSharePlugin_logic_mem_counter[3676] = 4'b0000;
    GSharePlugin_logic_mem_counter[3677] = 4'b0000;
    GSharePlugin_logic_mem_counter[3678] = 4'b0000;
    GSharePlugin_logic_mem_counter[3679] = 4'b0000;
    GSharePlugin_logic_mem_counter[3680] = 4'b0000;
    GSharePlugin_logic_mem_counter[3681] = 4'b0000;
    GSharePlugin_logic_mem_counter[3682] = 4'b0000;
    GSharePlugin_logic_mem_counter[3683] = 4'b0000;
    GSharePlugin_logic_mem_counter[3684] = 4'b0000;
    GSharePlugin_logic_mem_counter[3685] = 4'b0000;
    GSharePlugin_logic_mem_counter[3686] = 4'b0000;
    GSharePlugin_logic_mem_counter[3687] = 4'b0000;
    GSharePlugin_logic_mem_counter[3688] = 4'b0000;
    GSharePlugin_logic_mem_counter[3689] = 4'b0000;
    GSharePlugin_logic_mem_counter[3690] = 4'b0000;
    GSharePlugin_logic_mem_counter[3691] = 4'b0000;
    GSharePlugin_logic_mem_counter[3692] = 4'b0000;
    GSharePlugin_logic_mem_counter[3693] = 4'b0000;
    GSharePlugin_logic_mem_counter[3694] = 4'b0000;
    GSharePlugin_logic_mem_counter[3695] = 4'b0000;
    GSharePlugin_logic_mem_counter[3696] = 4'b0000;
    GSharePlugin_logic_mem_counter[3697] = 4'b0000;
    GSharePlugin_logic_mem_counter[3698] = 4'b0000;
    GSharePlugin_logic_mem_counter[3699] = 4'b0000;
    GSharePlugin_logic_mem_counter[3700] = 4'b0000;
    GSharePlugin_logic_mem_counter[3701] = 4'b0000;
    GSharePlugin_logic_mem_counter[3702] = 4'b0000;
    GSharePlugin_logic_mem_counter[3703] = 4'b0000;
    GSharePlugin_logic_mem_counter[3704] = 4'b0000;
    GSharePlugin_logic_mem_counter[3705] = 4'b0000;
    GSharePlugin_logic_mem_counter[3706] = 4'b0000;
    GSharePlugin_logic_mem_counter[3707] = 4'b0000;
    GSharePlugin_logic_mem_counter[3708] = 4'b0000;
    GSharePlugin_logic_mem_counter[3709] = 4'b0000;
    GSharePlugin_logic_mem_counter[3710] = 4'b0000;
    GSharePlugin_logic_mem_counter[3711] = 4'b0000;
    GSharePlugin_logic_mem_counter[3712] = 4'b0000;
    GSharePlugin_logic_mem_counter[3713] = 4'b0000;
    GSharePlugin_logic_mem_counter[3714] = 4'b0000;
    GSharePlugin_logic_mem_counter[3715] = 4'b0000;
    GSharePlugin_logic_mem_counter[3716] = 4'b0000;
    GSharePlugin_logic_mem_counter[3717] = 4'b0000;
    GSharePlugin_logic_mem_counter[3718] = 4'b0000;
    GSharePlugin_logic_mem_counter[3719] = 4'b0000;
    GSharePlugin_logic_mem_counter[3720] = 4'b0000;
    GSharePlugin_logic_mem_counter[3721] = 4'b0000;
    GSharePlugin_logic_mem_counter[3722] = 4'b0000;
    GSharePlugin_logic_mem_counter[3723] = 4'b0000;
    GSharePlugin_logic_mem_counter[3724] = 4'b0000;
    GSharePlugin_logic_mem_counter[3725] = 4'b0000;
    GSharePlugin_logic_mem_counter[3726] = 4'b0000;
    GSharePlugin_logic_mem_counter[3727] = 4'b0000;
    GSharePlugin_logic_mem_counter[3728] = 4'b0000;
    GSharePlugin_logic_mem_counter[3729] = 4'b0000;
    GSharePlugin_logic_mem_counter[3730] = 4'b0000;
    GSharePlugin_logic_mem_counter[3731] = 4'b0000;
    GSharePlugin_logic_mem_counter[3732] = 4'b0000;
    GSharePlugin_logic_mem_counter[3733] = 4'b0000;
    GSharePlugin_logic_mem_counter[3734] = 4'b0000;
    GSharePlugin_logic_mem_counter[3735] = 4'b0000;
    GSharePlugin_logic_mem_counter[3736] = 4'b0000;
    GSharePlugin_logic_mem_counter[3737] = 4'b0000;
    GSharePlugin_logic_mem_counter[3738] = 4'b0000;
    GSharePlugin_logic_mem_counter[3739] = 4'b0000;
    GSharePlugin_logic_mem_counter[3740] = 4'b0000;
    GSharePlugin_logic_mem_counter[3741] = 4'b0000;
    GSharePlugin_logic_mem_counter[3742] = 4'b0000;
    GSharePlugin_logic_mem_counter[3743] = 4'b0000;
    GSharePlugin_logic_mem_counter[3744] = 4'b0000;
    GSharePlugin_logic_mem_counter[3745] = 4'b0000;
    GSharePlugin_logic_mem_counter[3746] = 4'b0000;
    GSharePlugin_logic_mem_counter[3747] = 4'b0000;
    GSharePlugin_logic_mem_counter[3748] = 4'b0000;
    GSharePlugin_logic_mem_counter[3749] = 4'b0000;
    GSharePlugin_logic_mem_counter[3750] = 4'b0000;
    GSharePlugin_logic_mem_counter[3751] = 4'b0000;
    GSharePlugin_logic_mem_counter[3752] = 4'b0000;
    GSharePlugin_logic_mem_counter[3753] = 4'b0000;
    GSharePlugin_logic_mem_counter[3754] = 4'b0000;
    GSharePlugin_logic_mem_counter[3755] = 4'b0000;
    GSharePlugin_logic_mem_counter[3756] = 4'b0000;
    GSharePlugin_logic_mem_counter[3757] = 4'b0000;
    GSharePlugin_logic_mem_counter[3758] = 4'b0000;
    GSharePlugin_logic_mem_counter[3759] = 4'b0000;
    GSharePlugin_logic_mem_counter[3760] = 4'b0000;
    GSharePlugin_logic_mem_counter[3761] = 4'b0000;
    GSharePlugin_logic_mem_counter[3762] = 4'b0000;
    GSharePlugin_logic_mem_counter[3763] = 4'b0000;
    GSharePlugin_logic_mem_counter[3764] = 4'b0000;
    GSharePlugin_logic_mem_counter[3765] = 4'b0000;
    GSharePlugin_logic_mem_counter[3766] = 4'b0000;
    GSharePlugin_logic_mem_counter[3767] = 4'b0000;
    GSharePlugin_logic_mem_counter[3768] = 4'b0000;
    GSharePlugin_logic_mem_counter[3769] = 4'b0000;
    GSharePlugin_logic_mem_counter[3770] = 4'b0000;
    GSharePlugin_logic_mem_counter[3771] = 4'b0000;
    GSharePlugin_logic_mem_counter[3772] = 4'b0000;
    GSharePlugin_logic_mem_counter[3773] = 4'b0000;
    GSharePlugin_logic_mem_counter[3774] = 4'b0000;
    GSharePlugin_logic_mem_counter[3775] = 4'b0000;
    GSharePlugin_logic_mem_counter[3776] = 4'b0000;
    GSharePlugin_logic_mem_counter[3777] = 4'b0000;
    GSharePlugin_logic_mem_counter[3778] = 4'b0000;
    GSharePlugin_logic_mem_counter[3779] = 4'b0000;
    GSharePlugin_logic_mem_counter[3780] = 4'b0000;
    GSharePlugin_logic_mem_counter[3781] = 4'b0000;
    GSharePlugin_logic_mem_counter[3782] = 4'b0000;
    GSharePlugin_logic_mem_counter[3783] = 4'b0000;
    GSharePlugin_logic_mem_counter[3784] = 4'b0000;
    GSharePlugin_logic_mem_counter[3785] = 4'b0000;
    GSharePlugin_logic_mem_counter[3786] = 4'b0000;
    GSharePlugin_logic_mem_counter[3787] = 4'b0000;
    GSharePlugin_logic_mem_counter[3788] = 4'b0000;
    GSharePlugin_logic_mem_counter[3789] = 4'b0000;
    GSharePlugin_logic_mem_counter[3790] = 4'b0000;
    GSharePlugin_logic_mem_counter[3791] = 4'b0000;
    GSharePlugin_logic_mem_counter[3792] = 4'b0000;
    GSharePlugin_logic_mem_counter[3793] = 4'b0000;
    GSharePlugin_logic_mem_counter[3794] = 4'b0000;
    GSharePlugin_logic_mem_counter[3795] = 4'b0000;
    GSharePlugin_logic_mem_counter[3796] = 4'b0000;
    GSharePlugin_logic_mem_counter[3797] = 4'b0000;
    GSharePlugin_logic_mem_counter[3798] = 4'b0000;
    GSharePlugin_logic_mem_counter[3799] = 4'b0000;
    GSharePlugin_logic_mem_counter[3800] = 4'b0000;
    GSharePlugin_logic_mem_counter[3801] = 4'b0000;
    GSharePlugin_logic_mem_counter[3802] = 4'b0000;
    GSharePlugin_logic_mem_counter[3803] = 4'b0000;
    GSharePlugin_logic_mem_counter[3804] = 4'b0000;
    GSharePlugin_logic_mem_counter[3805] = 4'b0000;
    GSharePlugin_logic_mem_counter[3806] = 4'b0000;
    GSharePlugin_logic_mem_counter[3807] = 4'b0000;
    GSharePlugin_logic_mem_counter[3808] = 4'b0000;
    GSharePlugin_logic_mem_counter[3809] = 4'b0000;
    GSharePlugin_logic_mem_counter[3810] = 4'b0000;
    GSharePlugin_logic_mem_counter[3811] = 4'b0000;
    GSharePlugin_logic_mem_counter[3812] = 4'b0000;
    GSharePlugin_logic_mem_counter[3813] = 4'b0000;
    GSharePlugin_logic_mem_counter[3814] = 4'b0000;
    GSharePlugin_logic_mem_counter[3815] = 4'b0000;
    GSharePlugin_logic_mem_counter[3816] = 4'b0000;
    GSharePlugin_logic_mem_counter[3817] = 4'b0000;
    GSharePlugin_logic_mem_counter[3818] = 4'b0000;
    GSharePlugin_logic_mem_counter[3819] = 4'b0000;
    GSharePlugin_logic_mem_counter[3820] = 4'b0000;
    GSharePlugin_logic_mem_counter[3821] = 4'b0000;
    GSharePlugin_logic_mem_counter[3822] = 4'b0000;
    GSharePlugin_logic_mem_counter[3823] = 4'b0000;
    GSharePlugin_logic_mem_counter[3824] = 4'b0000;
    GSharePlugin_logic_mem_counter[3825] = 4'b0000;
    GSharePlugin_logic_mem_counter[3826] = 4'b0000;
    GSharePlugin_logic_mem_counter[3827] = 4'b0000;
    GSharePlugin_logic_mem_counter[3828] = 4'b0000;
    GSharePlugin_logic_mem_counter[3829] = 4'b0000;
    GSharePlugin_logic_mem_counter[3830] = 4'b0000;
    GSharePlugin_logic_mem_counter[3831] = 4'b0000;
    GSharePlugin_logic_mem_counter[3832] = 4'b0000;
    GSharePlugin_logic_mem_counter[3833] = 4'b0000;
    GSharePlugin_logic_mem_counter[3834] = 4'b0000;
    GSharePlugin_logic_mem_counter[3835] = 4'b0000;
    GSharePlugin_logic_mem_counter[3836] = 4'b0000;
    GSharePlugin_logic_mem_counter[3837] = 4'b0000;
    GSharePlugin_logic_mem_counter[3838] = 4'b0000;
    GSharePlugin_logic_mem_counter[3839] = 4'b0000;
    GSharePlugin_logic_mem_counter[3840] = 4'b0000;
    GSharePlugin_logic_mem_counter[3841] = 4'b0000;
    GSharePlugin_logic_mem_counter[3842] = 4'b0000;
    GSharePlugin_logic_mem_counter[3843] = 4'b0000;
    GSharePlugin_logic_mem_counter[3844] = 4'b0000;
    GSharePlugin_logic_mem_counter[3845] = 4'b0000;
    GSharePlugin_logic_mem_counter[3846] = 4'b0000;
    GSharePlugin_logic_mem_counter[3847] = 4'b0000;
    GSharePlugin_logic_mem_counter[3848] = 4'b0000;
    GSharePlugin_logic_mem_counter[3849] = 4'b0000;
    GSharePlugin_logic_mem_counter[3850] = 4'b0000;
    GSharePlugin_logic_mem_counter[3851] = 4'b0000;
    GSharePlugin_logic_mem_counter[3852] = 4'b0000;
    GSharePlugin_logic_mem_counter[3853] = 4'b0000;
    GSharePlugin_logic_mem_counter[3854] = 4'b0000;
    GSharePlugin_logic_mem_counter[3855] = 4'b0000;
    GSharePlugin_logic_mem_counter[3856] = 4'b0000;
    GSharePlugin_logic_mem_counter[3857] = 4'b0000;
    GSharePlugin_logic_mem_counter[3858] = 4'b0000;
    GSharePlugin_logic_mem_counter[3859] = 4'b0000;
    GSharePlugin_logic_mem_counter[3860] = 4'b0000;
    GSharePlugin_logic_mem_counter[3861] = 4'b0000;
    GSharePlugin_logic_mem_counter[3862] = 4'b0000;
    GSharePlugin_logic_mem_counter[3863] = 4'b0000;
    GSharePlugin_logic_mem_counter[3864] = 4'b0000;
    GSharePlugin_logic_mem_counter[3865] = 4'b0000;
    GSharePlugin_logic_mem_counter[3866] = 4'b0000;
    GSharePlugin_logic_mem_counter[3867] = 4'b0000;
    GSharePlugin_logic_mem_counter[3868] = 4'b0000;
    GSharePlugin_logic_mem_counter[3869] = 4'b0000;
    GSharePlugin_logic_mem_counter[3870] = 4'b0000;
    GSharePlugin_logic_mem_counter[3871] = 4'b0000;
    GSharePlugin_logic_mem_counter[3872] = 4'b0000;
    GSharePlugin_logic_mem_counter[3873] = 4'b0000;
    GSharePlugin_logic_mem_counter[3874] = 4'b0000;
    GSharePlugin_logic_mem_counter[3875] = 4'b0000;
    GSharePlugin_logic_mem_counter[3876] = 4'b0000;
    GSharePlugin_logic_mem_counter[3877] = 4'b0000;
    GSharePlugin_logic_mem_counter[3878] = 4'b0000;
    GSharePlugin_logic_mem_counter[3879] = 4'b0000;
    GSharePlugin_logic_mem_counter[3880] = 4'b0000;
    GSharePlugin_logic_mem_counter[3881] = 4'b0000;
    GSharePlugin_logic_mem_counter[3882] = 4'b0000;
    GSharePlugin_logic_mem_counter[3883] = 4'b0000;
    GSharePlugin_logic_mem_counter[3884] = 4'b0000;
    GSharePlugin_logic_mem_counter[3885] = 4'b0000;
    GSharePlugin_logic_mem_counter[3886] = 4'b0000;
    GSharePlugin_logic_mem_counter[3887] = 4'b0000;
    GSharePlugin_logic_mem_counter[3888] = 4'b0000;
    GSharePlugin_logic_mem_counter[3889] = 4'b0000;
    GSharePlugin_logic_mem_counter[3890] = 4'b0000;
    GSharePlugin_logic_mem_counter[3891] = 4'b0000;
    GSharePlugin_logic_mem_counter[3892] = 4'b0000;
    GSharePlugin_logic_mem_counter[3893] = 4'b0000;
    GSharePlugin_logic_mem_counter[3894] = 4'b0000;
    GSharePlugin_logic_mem_counter[3895] = 4'b0000;
    GSharePlugin_logic_mem_counter[3896] = 4'b0000;
    GSharePlugin_logic_mem_counter[3897] = 4'b0000;
    GSharePlugin_logic_mem_counter[3898] = 4'b0000;
    GSharePlugin_logic_mem_counter[3899] = 4'b0000;
    GSharePlugin_logic_mem_counter[3900] = 4'b0000;
    GSharePlugin_logic_mem_counter[3901] = 4'b0000;
    GSharePlugin_logic_mem_counter[3902] = 4'b0000;
    GSharePlugin_logic_mem_counter[3903] = 4'b0000;
    GSharePlugin_logic_mem_counter[3904] = 4'b0000;
    GSharePlugin_logic_mem_counter[3905] = 4'b0000;
    GSharePlugin_logic_mem_counter[3906] = 4'b0000;
    GSharePlugin_logic_mem_counter[3907] = 4'b0000;
    GSharePlugin_logic_mem_counter[3908] = 4'b0000;
    GSharePlugin_logic_mem_counter[3909] = 4'b0000;
    GSharePlugin_logic_mem_counter[3910] = 4'b0000;
    GSharePlugin_logic_mem_counter[3911] = 4'b0000;
    GSharePlugin_logic_mem_counter[3912] = 4'b0000;
    GSharePlugin_logic_mem_counter[3913] = 4'b0000;
    GSharePlugin_logic_mem_counter[3914] = 4'b0000;
    GSharePlugin_logic_mem_counter[3915] = 4'b0000;
    GSharePlugin_logic_mem_counter[3916] = 4'b0000;
    GSharePlugin_logic_mem_counter[3917] = 4'b0000;
    GSharePlugin_logic_mem_counter[3918] = 4'b0000;
    GSharePlugin_logic_mem_counter[3919] = 4'b0000;
    GSharePlugin_logic_mem_counter[3920] = 4'b0000;
    GSharePlugin_logic_mem_counter[3921] = 4'b0000;
    GSharePlugin_logic_mem_counter[3922] = 4'b0000;
    GSharePlugin_logic_mem_counter[3923] = 4'b0000;
    GSharePlugin_logic_mem_counter[3924] = 4'b0000;
    GSharePlugin_logic_mem_counter[3925] = 4'b0000;
    GSharePlugin_logic_mem_counter[3926] = 4'b0000;
    GSharePlugin_logic_mem_counter[3927] = 4'b0000;
    GSharePlugin_logic_mem_counter[3928] = 4'b0000;
    GSharePlugin_logic_mem_counter[3929] = 4'b0000;
    GSharePlugin_logic_mem_counter[3930] = 4'b0000;
    GSharePlugin_logic_mem_counter[3931] = 4'b0000;
    GSharePlugin_logic_mem_counter[3932] = 4'b0000;
    GSharePlugin_logic_mem_counter[3933] = 4'b0000;
    GSharePlugin_logic_mem_counter[3934] = 4'b0000;
    GSharePlugin_logic_mem_counter[3935] = 4'b0000;
    GSharePlugin_logic_mem_counter[3936] = 4'b0000;
    GSharePlugin_logic_mem_counter[3937] = 4'b0000;
    GSharePlugin_logic_mem_counter[3938] = 4'b0000;
    GSharePlugin_logic_mem_counter[3939] = 4'b0000;
    GSharePlugin_logic_mem_counter[3940] = 4'b0000;
    GSharePlugin_logic_mem_counter[3941] = 4'b0000;
    GSharePlugin_logic_mem_counter[3942] = 4'b0000;
    GSharePlugin_logic_mem_counter[3943] = 4'b0000;
    GSharePlugin_logic_mem_counter[3944] = 4'b0000;
    GSharePlugin_logic_mem_counter[3945] = 4'b0000;
    GSharePlugin_logic_mem_counter[3946] = 4'b0000;
    GSharePlugin_logic_mem_counter[3947] = 4'b0000;
    GSharePlugin_logic_mem_counter[3948] = 4'b0000;
    GSharePlugin_logic_mem_counter[3949] = 4'b0000;
    GSharePlugin_logic_mem_counter[3950] = 4'b0000;
    GSharePlugin_logic_mem_counter[3951] = 4'b0000;
    GSharePlugin_logic_mem_counter[3952] = 4'b0000;
    GSharePlugin_logic_mem_counter[3953] = 4'b0000;
    GSharePlugin_logic_mem_counter[3954] = 4'b0000;
    GSharePlugin_logic_mem_counter[3955] = 4'b0000;
    GSharePlugin_logic_mem_counter[3956] = 4'b0000;
    GSharePlugin_logic_mem_counter[3957] = 4'b0000;
    GSharePlugin_logic_mem_counter[3958] = 4'b0000;
    GSharePlugin_logic_mem_counter[3959] = 4'b0000;
    GSharePlugin_logic_mem_counter[3960] = 4'b0000;
    GSharePlugin_logic_mem_counter[3961] = 4'b0000;
    GSharePlugin_logic_mem_counter[3962] = 4'b0000;
    GSharePlugin_logic_mem_counter[3963] = 4'b0000;
    GSharePlugin_logic_mem_counter[3964] = 4'b0000;
    GSharePlugin_logic_mem_counter[3965] = 4'b0000;
    GSharePlugin_logic_mem_counter[3966] = 4'b0000;
    GSharePlugin_logic_mem_counter[3967] = 4'b0000;
    GSharePlugin_logic_mem_counter[3968] = 4'b0000;
    GSharePlugin_logic_mem_counter[3969] = 4'b0000;
    GSharePlugin_logic_mem_counter[3970] = 4'b0000;
    GSharePlugin_logic_mem_counter[3971] = 4'b0000;
    GSharePlugin_logic_mem_counter[3972] = 4'b0000;
    GSharePlugin_logic_mem_counter[3973] = 4'b0000;
    GSharePlugin_logic_mem_counter[3974] = 4'b0000;
    GSharePlugin_logic_mem_counter[3975] = 4'b0000;
    GSharePlugin_logic_mem_counter[3976] = 4'b0000;
    GSharePlugin_logic_mem_counter[3977] = 4'b0000;
    GSharePlugin_logic_mem_counter[3978] = 4'b0000;
    GSharePlugin_logic_mem_counter[3979] = 4'b0000;
    GSharePlugin_logic_mem_counter[3980] = 4'b0000;
    GSharePlugin_logic_mem_counter[3981] = 4'b0000;
    GSharePlugin_logic_mem_counter[3982] = 4'b0000;
    GSharePlugin_logic_mem_counter[3983] = 4'b0000;
    GSharePlugin_logic_mem_counter[3984] = 4'b0000;
    GSharePlugin_logic_mem_counter[3985] = 4'b0000;
    GSharePlugin_logic_mem_counter[3986] = 4'b0000;
    GSharePlugin_logic_mem_counter[3987] = 4'b0000;
    GSharePlugin_logic_mem_counter[3988] = 4'b0000;
    GSharePlugin_logic_mem_counter[3989] = 4'b0000;
    GSharePlugin_logic_mem_counter[3990] = 4'b0000;
    GSharePlugin_logic_mem_counter[3991] = 4'b0000;
    GSharePlugin_logic_mem_counter[3992] = 4'b0000;
    GSharePlugin_logic_mem_counter[3993] = 4'b0000;
    GSharePlugin_logic_mem_counter[3994] = 4'b0000;
    GSharePlugin_logic_mem_counter[3995] = 4'b0000;
    GSharePlugin_logic_mem_counter[3996] = 4'b0000;
    GSharePlugin_logic_mem_counter[3997] = 4'b0000;
    GSharePlugin_logic_mem_counter[3998] = 4'b0000;
    GSharePlugin_logic_mem_counter[3999] = 4'b0000;
    GSharePlugin_logic_mem_counter[4000] = 4'b0000;
    GSharePlugin_logic_mem_counter[4001] = 4'b0000;
    GSharePlugin_logic_mem_counter[4002] = 4'b0000;
    GSharePlugin_logic_mem_counter[4003] = 4'b0000;
    GSharePlugin_logic_mem_counter[4004] = 4'b0000;
    GSharePlugin_logic_mem_counter[4005] = 4'b0000;
    GSharePlugin_logic_mem_counter[4006] = 4'b0000;
    GSharePlugin_logic_mem_counter[4007] = 4'b0000;
    GSharePlugin_logic_mem_counter[4008] = 4'b0000;
    GSharePlugin_logic_mem_counter[4009] = 4'b0000;
    GSharePlugin_logic_mem_counter[4010] = 4'b0000;
    GSharePlugin_logic_mem_counter[4011] = 4'b0000;
    GSharePlugin_logic_mem_counter[4012] = 4'b0000;
    GSharePlugin_logic_mem_counter[4013] = 4'b0000;
    GSharePlugin_logic_mem_counter[4014] = 4'b0000;
    GSharePlugin_logic_mem_counter[4015] = 4'b0000;
    GSharePlugin_logic_mem_counter[4016] = 4'b0000;
    GSharePlugin_logic_mem_counter[4017] = 4'b0000;
    GSharePlugin_logic_mem_counter[4018] = 4'b0000;
    GSharePlugin_logic_mem_counter[4019] = 4'b0000;
    GSharePlugin_logic_mem_counter[4020] = 4'b0000;
    GSharePlugin_logic_mem_counter[4021] = 4'b0000;
    GSharePlugin_logic_mem_counter[4022] = 4'b0000;
    GSharePlugin_logic_mem_counter[4023] = 4'b0000;
    GSharePlugin_logic_mem_counter[4024] = 4'b0000;
    GSharePlugin_logic_mem_counter[4025] = 4'b0000;
    GSharePlugin_logic_mem_counter[4026] = 4'b0000;
    GSharePlugin_logic_mem_counter[4027] = 4'b0000;
    GSharePlugin_logic_mem_counter[4028] = 4'b0000;
    GSharePlugin_logic_mem_counter[4029] = 4'b0000;
    GSharePlugin_logic_mem_counter[4030] = 4'b0000;
    GSharePlugin_logic_mem_counter[4031] = 4'b0000;
    GSharePlugin_logic_mem_counter[4032] = 4'b0000;
    GSharePlugin_logic_mem_counter[4033] = 4'b0000;
    GSharePlugin_logic_mem_counter[4034] = 4'b0000;
    GSharePlugin_logic_mem_counter[4035] = 4'b0000;
    GSharePlugin_logic_mem_counter[4036] = 4'b0000;
    GSharePlugin_logic_mem_counter[4037] = 4'b0000;
    GSharePlugin_logic_mem_counter[4038] = 4'b0000;
    GSharePlugin_logic_mem_counter[4039] = 4'b0000;
    GSharePlugin_logic_mem_counter[4040] = 4'b0000;
    GSharePlugin_logic_mem_counter[4041] = 4'b0000;
    GSharePlugin_logic_mem_counter[4042] = 4'b0000;
    GSharePlugin_logic_mem_counter[4043] = 4'b0000;
    GSharePlugin_logic_mem_counter[4044] = 4'b0000;
    GSharePlugin_logic_mem_counter[4045] = 4'b0000;
    GSharePlugin_logic_mem_counter[4046] = 4'b0000;
    GSharePlugin_logic_mem_counter[4047] = 4'b0000;
    GSharePlugin_logic_mem_counter[4048] = 4'b0000;
    GSharePlugin_logic_mem_counter[4049] = 4'b0000;
    GSharePlugin_logic_mem_counter[4050] = 4'b0000;
    GSharePlugin_logic_mem_counter[4051] = 4'b0000;
    GSharePlugin_logic_mem_counter[4052] = 4'b0000;
    GSharePlugin_logic_mem_counter[4053] = 4'b0000;
    GSharePlugin_logic_mem_counter[4054] = 4'b0000;
    GSharePlugin_logic_mem_counter[4055] = 4'b0000;
    GSharePlugin_logic_mem_counter[4056] = 4'b0000;
    GSharePlugin_logic_mem_counter[4057] = 4'b0000;
    GSharePlugin_logic_mem_counter[4058] = 4'b0000;
    GSharePlugin_logic_mem_counter[4059] = 4'b0000;
    GSharePlugin_logic_mem_counter[4060] = 4'b0000;
    GSharePlugin_logic_mem_counter[4061] = 4'b0000;
    GSharePlugin_logic_mem_counter[4062] = 4'b0000;
    GSharePlugin_logic_mem_counter[4063] = 4'b0000;
    GSharePlugin_logic_mem_counter[4064] = 4'b0000;
    GSharePlugin_logic_mem_counter[4065] = 4'b0000;
    GSharePlugin_logic_mem_counter[4066] = 4'b0000;
    GSharePlugin_logic_mem_counter[4067] = 4'b0000;
    GSharePlugin_logic_mem_counter[4068] = 4'b0000;
    GSharePlugin_logic_mem_counter[4069] = 4'b0000;
    GSharePlugin_logic_mem_counter[4070] = 4'b0000;
    GSharePlugin_logic_mem_counter[4071] = 4'b0000;
    GSharePlugin_logic_mem_counter[4072] = 4'b0000;
    GSharePlugin_logic_mem_counter[4073] = 4'b0000;
    GSharePlugin_logic_mem_counter[4074] = 4'b0000;
    GSharePlugin_logic_mem_counter[4075] = 4'b0000;
    GSharePlugin_logic_mem_counter[4076] = 4'b0000;
    GSharePlugin_logic_mem_counter[4077] = 4'b0000;
    GSharePlugin_logic_mem_counter[4078] = 4'b0000;
    GSharePlugin_logic_mem_counter[4079] = 4'b0000;
    GSharePlugin_logic_mem_counter[4080] = 4'b0000;
    GSharePlugin_logic_mem_counter[4081] = 4'b0000;
    GSharePlugin_logic_mem_counter[4082] = 4'b0000;
    GSharePlugin_logic_mem_counter[4083] = 4'b0000;
    GSharePlugin_logic_mem_counter[4084] = 4'b0000;
    GSharePlugin_logic_mem_counter[4085] = 4'b0000;
    GSharePlugin_logic_mem_counter[4086] = 4'b0000;
    GSharePlugin_logic_mem_counter[4087] = 4'b0000;
    GSharePlugin_logic_mem_counter[4088] = 4'b0000;
    GSharePlugin_logic_mem_counter[4089] = 4'b0000;
    GSharePlugin_logic_mem_counter[4090] = 4'b0000;
    GSharePlugin_logic_mem_counter[4091] = 4'b0000;
    GSharePlugin_logic_mem_counter[4092] = 4'b0000;
    GSharePlugin_logic_mem_counter[4093] = 4'b0000;
    GSharePlugin_logic_mem_counter[4094] = 4'b0000;
    GSharePlugin_logic_mem_counter[4095] = 4'b0000;
    GSharePlugin_logic_mem_counter[4096] = 4'b0000;
    GSharePlugin_logic_mem_counter[4097] = 4'b0000;
    GSharePlugin_logic_mem_counter[4098] = 4'b0000;
    GSharePlugin_logic_mem_counter[4099] = 4'b0000;
    GSharePlugin_logic_mem_counter[4100] = 4'b0000;
    GSharePlugin_logic_mem_counter[4101] = 4'b0000;
    GSharePlugin_logic_mem_counter[4102] = 4'b0000;
    GSharePlugin_logic_mem_counter[4103] = 4'b0000;
    GSharePlugin_logic_mem_counter[4104] = 4'b0000;
    GSharePlugin_logic_mem_counter[4105] = 4'b0000;
    GSharePlugin_logic_mem_counter[4106] = 4'b0000;
    GSharePlugin_logic_mem_counter[4107] = 4'b0000;
    GSharePlugin_logic_mem_counter[4108] = 4'b0000;
    GSharePlugin_logic_mem_counter[4109] = 4'b0000;
    GSharePlugin_logic_mem_counter[4110] = 4'b0000;
    GSharePlugin_logic_mem_counter[4111] = 4'b0000;
    GSharePlugin_logic_mem_counter[4112] = 4'b0000;
    GSharePlugin_logic_mem_counter[4113] = 4'b0000;
    GSharePlugin_logic_mem_counter[4114] = 4'b0000;
    GSharePlugin_logic_mem_counter[4115] = 4'b0000;
    GSharePlugin_logic_mem_counter[4116] = 4'b0000;
    GSharePlugin_logic_mem_counter[4117] = 4'b0000;
    GSharePlugin_logic_mem_counter[4118] = 4'b0000;
    GSharePlugin_logic_mem_counter[4119] = 4'b0000;
    GSharePlugin_logic_mem_counter[4120] = 4'b0000;
    GSharePlugin_logic_mem_counter[4121] = 4'b0000;
    GSharePlugin_logic_mem_counter[4122] = 4'b0000;
    GSharePlugin_logic_mem_counter[4123] = 4'b0000;
    GSharePlugin_logic_mem_counter[4124] = 4'b0000;
    GSharePlugin_logic_mem_counter[4125] = 4'b0000;
    GSharePlugin_logic_mem_counter[4126] = 4'b0000;
    GSharePlugin_logic_mem_counter[4127] = 4'b0000;
    GSharePlugin_logic_mem_counter[4128] = 4'b0000;
    GSharePlugin_logic_mem_counter[4129] = 4'b0000;
    GSharePlugin_logic_mem_counter[4130] = 4'b0000;
    GSharePlugin_logic_mem_counter[4131] = 4'b0000;
    GSharePlugin_logic_mem_counter[4132] = 4'b0000;
    GSharePlugin_logic_mem_counter[4133] = 4'b0000;
    GSharePlugin_logic_mem_counter[4134] = 4'b0000;
    GSharePlugin_logic_mem_counter[4135] = 4'b0000;
    GSharePlugin_logic_mem_counter[4136] = 4'b0000;
    GSharePlugin_logic_mem_counter[4137] = 4'b0000;
    GSharePlugin_logic_mem_counter[4138] = 4'b0000;
    GSharePlugin_logic_mem_counter[4139] = 4'b0000;
    GSharePlugin_logic_mem_counter[4140] = 4'b0000;
    GSharePlugin_logic_mem_counter[4141] = 4'b0000;
    GSharePlugin_logic_mem_counter[4142] = 4'b0000;
    GSharePlugin_logic_mem_counter[4143] = 4'b0000;
    GSharePlugin_logic_mem_counter[4144] = 4'b0000;
    GSharePlugin_logic_mem_counter[4145] = 4'b0000;
    GSharePlugin_logic_mem_counter[4146] = 4'b0000;
    GSharePlugin_logic_mem_counter[4147] = 4'b0000;
    GSharePlugin_logic_mem_counter[4148] = 4'b0000;
    GSharePlugin_logic_mem_counter[4149] = 4'b0000;
    GSharePlugin_logic_mem_counter[4150] = 4'b0000;
    GSharePlugin_logic_mem_counter[4151] = 4'b0000;
    GSharePlugin_logic_mem_counter[4152] = 4'b0000;
    GSharePlugin_logic_mem_counter[4153] = 4'b0000;
    GSharePlugin_logic_mem_counter[4154] = 4'b0000;
    GSharePlugin_logic_mem_counter[4155] = 4'b0000;
    GSharePlugin_logic_mem_counter[4156] = 4'b0000;
    GSharePlugin_logic_mem_counter[4157] = 4'b0000;
    GSharePlugin_logic_mem_counter[4158] = 4'b0000;
    GSharePlugin_logic_mem_counter[4159] = 4'b0000;
    GSharePlugin_logic_mem_counter[4160] = 4'b0000;
    GSharePlugin_logic_mem_counter[4161] = 4'b0000;
    GSharePlugin_logic_mem_counter[4162] = 4'b0000;
    GSharePlugin_logic_mem_counter[4163] = 4'b0000;
    GSharePlugin_logic_mem_counter[4164] = 4'b0000;
    GSharePlugin_logic_mem_counter[4165] = 4'b0000;
    GSharePlugin_logic_mem_counter[4166] = 4'b0000;
    GSharePlugin_logic_mem_counter[4167] = 4'b0000;
    GSharePlugin_logic_mem_counter[4168] = 4'b0000;
    GSharePlugin_logic_mem_counter[4169] = 4'b0000;
    GSharePlugin_logic_mem_counter[4170] = 4'b0000;
    GSharePlugin_logic_mem_counter[4171] = 4'b0000;
    GSharePlugin_logic_mem_counter[4172] = 4'b0000;
    GSharePlugin_logic_mem_counter[4173] = 4'b0000;
    GSharePlugin_logic_mem_counter[4174] = 4'b0000;
    GSharePlugin_logic_mem_counter[4175] = 4'b0000;
    GSharePlugin_logic_mem_counter[4176] = 4'b0000;
    GSharePlugin_logic_mem_counter[4177] = 4'b0000;
    GSharePlugin_logic_mem_counter[4178] = 4'b0000;
    GSharePlugin_logic_mem_counter[4179] = 4'b0000;
    GSharePlugin_logic_mem_counter[4180] = 4'b0000;
    GSharePlugin_logic_mem_counter[4181] = 4'b0000;
    GSharePlugin_logic_mem_counter[4182] = 4'b0000;
    GSharePlugin_logic_mem_counter[4183] = 4'b0000;
    GSharePlugin_logic_mem_counter[4184] = 4'b0000;
    GSharePlugin_logic_mem_counter[4185] = 4'b0000;
    GSharePlugin_logic_mem_counter[4186] = 4'b0000;
    GSharePlugin_logic_mem_counter[4187] = 4'b0000;
    GSharePlugin_logic_mem_counter[4188] = 4'b0000;
    GSharePlugin_logic_mem_counter[4189] = 4'b0000;
    GSharePlugin_logic_mem_counter[4190] = 4'b0000;
    GSharePlugin_logic_mem_counter[4191] = 4'b0000;
    GSharePlugin_logic_mem_counter[4192] = 4'b0000;
    GSharePlugin_logic_mem_counter[4193] = 4'b0000;
    GSharePlugin_logic_mem_counter[4194] = 4'b0000;
    GSharePlugin_logic_mem_counter[4195] = 4'b0000;
    GSharePlugin_logic_mem_counter[4196] = 4'b0000;
    GSharePlugin_logic_mem_counter[4197] = 4'b0000;
    GSharePlugin_logic_mem_counter[4198] = 4'b0000;
    GSharePlugin_logic_mem_counter[4199] = 4'b0000;
    GSharePlugin_logic_mem_counter[4200] = 4'b0000;
    GSharePlugin_logic_mem_counter[4201] = 4'b0000;
    GSharePlugin_logic_mem_counter[4202] = 4'b0000;
    GSharePlugin_logic_mem_counter[4203] = 4'b0000;
    GSharePlugin_logic_mem_counter[4204] = 4'b0000;
    GSharePlugin_logic_mem_counter[4205] = 4'b0000;
    GSharePlugin_logic_mem_counter[4206] = 4'b0000;
    GSharePlugin_logic_mem_counter[4207] = 4'b0000;
    GSharePlugin_logic_mem_counter[4208] = 4'b0000;
    GSharePlugin_logic_mem_counter[4209] = 4'b0000;
    GSharePlugin_logic_mem_counter[4210] = 4'b0000;
    GSharePlugin_logic_mem_counter[4211] = 4'b0000;
    GSharePlugin_logic_mem_counter[4212] = 4'b0000;
    GSharePlugin_logic_mem_counter[4213] = 4'b0000;
    GSharePlugin_logic_mem_counter[4214] = 4'b0000;
    GSharePlugin_logic_mem_counter[4215] = 4'b0000;
    GSharePlugin_logic_mem_counter[4216] = 4'b0000;
    GSharePlugin_logic_mem_counter[4217] = 4'b0000;
    GSharePlugin_logic_mem_counter[4218] = 4'b0000;
    GSharePlugin_logic_mem_counter[4219] = 4'b0000;
    GSharePlugin_logic_mem_counter[4220] = 4'b0000;
    GSharePlugin_logic_mem_counter[4221] = 4'b0000;
    GSharePlugin_logic_mem_counter[4222] = 4'b0000;
    GSharePlugin_logic_mem_counter[4223] = 4'b0000;
    GSharePlugin_logic_mem_counter[4224] = 4'b0000;
    GSharePlugin_logic_mem_counter[4225] = 4'b0000;
    GSharePlugin_logic_mem_counter[4226] = 4'b0000;
    GSharePlugin_logic_mem_counter[4227] = 4'b0000;
    GSharePlugin_logic_mem_counter[4228] = 4'b0000;
    GSharePlugin_logic_mem_counter[4229] = 4'b0000;
    GSharePlugin_logic_mem_counter[4230] = 4'b0000;
    GSharePlugin_logic_mem_counter[4231] = 4'b0000;
    GSharePlugin_logic_mem_counter[4232] = 4'b0000;
    GSharePlugin_logic_mem_counter[4233] = 4'b0000;
    GSharePlugin_logic_mem_counter[4234] = 4'b0000;
    GSharePlugin_logic_mem_counter[4235] = 4'b0000;
    GSharePlugin_logic_mem_counter[4236] = 4'b0000;
    GSharePlugin_logic_mem_counter[4237] = 4'b0000;
    GSharePlugin_logic_mem_counter[4238] = 4'b0000;
    GSharePlugin_logic_mem_counter[4239] = 4'b0000;
    GSharePlugin_logic_mem_counter[4240] = 4'b0000;
    GSharePlugin_logic_mem_counter[4241] = 4'b0000;
    GSharePlugin_logic_mem_counter[4242] = 4'b0000;
    GSharePlugin_logic_mem_counter[4243] = 4'b0000;
    GSharePlugin_logic_mem_counter[4244] = 4'b0000;
    GSharePlugin_logic_mem_counter[4245] = 4'b0000;
    GSharePlugin_logic_mem_counter[4246] = 4'b0000;
    GSharePlugin_logic_mem_counter[4247] = 4'b0000;
    GSharePlugin_logic_mem_counter[4248] = 4'b0000;
    GSharePlugin_logic_mem_counter[4249] = 4'b0000;
    GSharePlugin_logic_mem_counter[4250] = 4'b0000;
    GSharePlugin_logic_mem_counter[4251] = 4'b0000;
    GSharePlugin_logic_mem_counter[4252] = 4'b0000;
    GSharePlugin_logic_mem_counter[4253] = 4'b0000;
    GSharePlugin_logic_mem_counter[4254] = 4'b0000;
    GSharePlugin_logic_mem_counter[4255] = 4'b0000;
    GSharePlugin_logic_mem_counter[4256] = 4'b0000;
    GSharePlugin_logic_mem_counter[4257] = 4'b0000;
    GSharePlugin_logic_mem_counter[4258] = 4'b0000;
    GSharePlugin_logic_mem_counter[4259] = 4'b0000;
    GSharePlugin_logic_mem_counter[4260] = 4'b0000;
    GSharePlugin_logic_mem_counter[4261] = 4'b0000;
    GSharePlugin_logic_mem_counter[4262] = 4'b0000;
    GSharePlugin_logic_mem_counter[4263] = 4'b0000;
    GSharePlugin_logic_mem_counter[4264] = 4'b0000;
    GSharePlugin_logic_mem_counter[4265] = 4'b0000;
    GSharePlugin_logic_mem_counter[4266] = 4'b0000;
    GSharePlugin_logic_mem_counter[4267] = 4'b0000;
    GSharePlugin_logic_mem_counter[4268] = 4'b0000;
    GSharePlugin_logic_mem_counter[4269] = 4'b0000;
    GSharePlugin_logic_mem_counter[4270] = 4'b0000;
    GSharePlugin_logic_mem_counter[4271] = 4'b0000;
    GSharePlugin_logic_mem_counter[4272] = 4'b0000;
    GSharePlugin_logic_mem_counter[4273] = 4'b0000;
    GSharePlugin_logic_mem_counter[4274] = 4'b0000;
    GSharePlugin_logic_mem_counter[4275] = 4'b0000;
    GSharePlugin_logic_mem_counter[4276] = 4'b0000;
    GSharePlugin_logic_mem_counter[4277] = 4'b0000;
    GSharePlugin_logic_mem_counter[4278] = 4'b0000;
    GSharePlugin_logic_mem_counter[4279] = 4'b0000;
    GSharePlugin_logic_mem_counter[4280] = 4'b0000;
    GSharePlugin_logic_mem_counter[4281] = 4'b0000;
    GSharePlugin_logic_mem_counter[4282] = 4'b0000;
    GSharePlugin_logic_mem_counter[4283] = 4'b0000;
    GSharePlugin_logic_mem_counter[4284] = 4'b0000;
    GSharePlugin_logic_mem_counter[4285] = 4'b0000;
    GSharePlugin_logic_mem_counter[4286] = 4'b0000;
    GSharePlugin_logic_mem_counter[4287] = 4'b0000;
    GSharePlugin_logic_mem_counter[4288] = 4'b0000;
    GSharePlugin_logic_mem_counter[4289] = 4'b0000;
    GSharePlugin_logic_mem_counter[4290] = 4'b0000;
    GSharePlugin_logic_mem_counter[4291] = 4'b0000;
    GSharePlugin_logic_mem_counter[4292] = 4'b0000;
    GSharePlugin_logic_mem_counter[4293] = 4'b0000;
    GSharePlugin_logic_mem_counter[4294] = 4'b0000;
    GSharePlugin_logic_mem_counter[4295] = 4'b0000;
    GSharePlugin_logic_mem_counter[4296] = 4'b0000;
    GSharePlugin_logic_mem_counter[4297] = 4'b0000;
    GSharePlugin_logic_mem_counter[4298] = 4'b0000;
    GSharePlugin_logic_mem_counter[4299] = 4'b0000;
    GSharePlugin_logic_mem_counter[4300] = 4'b0000;
    GSharePlugin_logic_mem_counter[4301] = 4'b0000;
    GSharePlugin_logic_mem_counter[4302] = 4'b0000;
    GSharePlugin_logic_mem_counter[4303] = 4'b0000;
    GSharePlugin_logic_mem_counter[4304] = 4'b0000;
    GSharePlugin_logic_mem_counter[4305] = 4'b0000;
    GSharePlugin_logic_mem_counter[4306] = 4'b0000;
    GSharePlugin_logic_mem_counter[4307] = 4'b0000;
    GSharePlugin_logic_mem_counter[4308] = 4'b0000;
    GSharePlugin_logic_mem_counter[4309] = 4'b0000;
    GSharePlugin_logic_mem_counter[4310] = 4'b0000;
    GSharePlugin_logic_mem_counter[4311] = 4'b0000;
    GSharePlugin_logic_mem_counter[4312] = 4'b0000;
    GSharePlugin_logic_mem_counter[4313] = 4'b0000;
    GSharePlugin_logic_mem_counter[4314] = 4'b0000;
    GSharePlugin_logic_mem_counter[4315] = 4'b0000;
    GSharePlugin_logic_mem_counter[4316] = 4'b0000;
    GSharePlugin_logic_mem_counter[4317] = 4'b0000;
    GSharePlugin_logic_mem_counter[4318] = 4'b0000;
    GSharePlugin_logic_mem_counter[4319] = 4'b0000;
    GSharePlugin_logic_mem_counter[4320] = 4'b0000;
    GSharePlugin_logic_mem_counter[4321] = 4'b0000;
    GSharePlugin_logic_mem_counter[4322] = 4'b0000;
    GSharePlugin_logic_mem_counter[4323] = 4'b0000;
    GSharePlugin_logic_mem_counter[4324] = 4'b0000;
    GSharePlugin_logic_mem_counter[4325] = 4'b0000;
    GSharePlugin_logic_mem_counter[4326] = 4'b0000;
    GSharePlugin_logic_mem_counter[4327] = 4'b0000;
    GSharePlugin_logic_mem_counter[4328] = 4'b0000;
    GSharePlugin_logic_mem_counter[4329] = 4'b0000;
    GSharePlugin_logic_mem_counter[4330] = 4'b0000;
    GSharePlugin_logic_mem_counter[4331] = 4'b0000;
    GSharePlugin_logic_mem_counter[4332] = 4'b0000;
    GSharePlugin_logic_mem_counter[4333] = 4'b0000;
    GSharePlugin_logic_mem_counter[4334] = 4'b0000;
    GSharePlugin_logic_mem_counter[4335] = 4'b0000;
    GSharePlugin_logic_mem_counter[4336] = 4'b0000;
    GSharePlugin_logic_mem_counter[4337] = 4'b0000;
    GSharePlugin_logic_mem_counter[4338] = 4'b0000;
    GSharePlugin_logic_mem_counter[4339] = 4'b0000;
    GSharePlugin_logic_mem_counter[4340] = 4'b0000;
    GSharePlugin_logic_mem_counter[4341] = 4'b0000;
    GSharePlugin_logic_mem_counter[4342] = 4'b0000;
    GSharePlugin_logic_mem_counter[4343] = 4'b0000;
    GSharePlugin_logic_mem_counter[4344] = 4'b0000;
    GSharePlugin_logic_mem_counter[4345] = 4'b0000;
    GSharePlugin_logic_mem_counter[4346] = 4'b0000;
    GSharePlugin_logic_mem_counter[4347] = 4'b0000;
    GSharePlugin_logic_mem_counter[4348] = 4'b0000;
    GSharePlugin_logic_mem_counter[4349] = 4'b0000;
    GSharePlugin_logic_mem_counter[4350] = 4'b0000;
    GSharePlugin_logic_mem_counter[4351] = 4'b0000;
    GSharePlugin_logic_mem_counter[4352] = 4'b0000;
    GSharePlugin_logic_mem_counter[4353] = 4'b0000;
    GSharePlugin_logic_mem_counter[4354] = 4'b0000;
    GSharePlugin_logic_mem_counter[4355] = 4'b0000;
    GSharePlugin_logic_mem_counter[4356] = 4'b0000;
    GSharePlugin_logic_mem_counter[4357] = 4'b0000;
    GSharePlugin_logic_mem_counter[4358] = 4'b0000;
    GSharePlugin_logic_mem_counter[4359] = 4'b0000;
    GSharePlugin_logic_mem_counter[4360] = 4'b0000;
    GSharePlugin_logic_mem_counter[4361] = 4'b0000;
    GSharePlugin_logic_mem_counter[4362] = 4'b0000;
    GSharePlugin_logic_mem_counter[4363] = 4'b0000;
    GSharePlugin_logic_mem_counter[4364] = 4'b0000;
    GSharePlugin_logic_mem_counter[4365] = 4'b0000;
    GSharePlugin_logic_mem_counter[4366] = 4'b0000;
    GSharePlugin_logic_mem_counter[4367] = 4'b0000;
    GSharePlugin_logic_mem_counter[4368] = 4'b0000;
    GSharePlugin_logic_mem_counter[4369] = 4'b0000;
    GSharePlugin_logic_mem_counter[4370] = 4'b0000;
    GSharePlugin_logic_mem_counter[4371] = 4'b0000;
    GSharePlugin_logic_mem_counter[4372] = 4'b0000;
    GSharePlugin_logic_mem_counter[4373] = 4'b0000;
    GSharePlugin_logic_mem_counter[4374] = 4'b0000;
    GSharePlugin_logic_mem_counter[4375] = 4'b0000;
    GSharePlugin_logic_mem_counter[4376] = 4'b0000;
    GSharePlugin_logic_mem_counter[4377] = 4'b0000;
    GSharePlugin_logic_mem_counter[4378] = 4'b0000;
    GSharePlugin_logic_mem_counter[4379] = 4'b0000;
    GSharePlugin_logic_mem_counter[4380] = 4'b0000;
    GSharePlugin_logic_mem_counter[4381] = 4'b0000;
    GSharePlugin_logic_mem_counter[4382] = 4'b0000;
    GSharePlugin_logic_mem_counter[4383] = 4'b0000;
    GSharePlugin_logic_mem_counter[4384] = 4'b0000;
    GSharePlugin_logic_mem_counter[4385] = 4'b0000;
    GSharePlugin_logic_mem_counter[4386] = 4'b0000;
    GSharePlugin_logic_mem_counter[4387] = 4'b0000;
    GSharePlugin_logic_mem_counter[4388] = 4'b0000;
    GSharePlugin_logic_mem_counter[4389] = 4'b0000;
    GSharePlugin_logic_mem_counter[4390] = 4'b0000;
    GSharePlugin_logic_mem_counter[4391] = 4'b0000;
    GSharePlugin_logic_mem_counter[4392] = 4'b0000;
    GSharePlugin_logic_mem_counter[4393] = 4'b0000;
    GSharePlugin_logic_mem_counter[4394] = 4'b0000;
    GSharePlugin_logic_mem_counter[4395] = 4'b0000;
    GSharePlugin_logic_mem_counter[4396] = 4'b0000;
    GSharePlugin_logic_mem_counter[4397] = 4'b0000;
    GSharePlugin_logic_mem_counter[4398] = 4'b0000;
    GSharePlugin_logic_mem_counter[4399] = 4'b0000;
    GSharePlugin_logic_mem_counter[4400] = 4'b0000;
    GSharePlugin_logic_mem_counter[4401] = 4'b0000;
    GSharePlugin_logic_mem_counter[4402] = 4'b0000;
    GSharePlugin_logic_mem_counter[4403] = 4'b0000;
    GSharePlugin_logic_mem_counter[4404] = 4'b0000;
    GSharePlugin_logic_mem_counter[4405] = 4'b0000;
    GSharePlugin_logic_mem_counter[4406] = 4'b0000;
    GSharePlugin_logic_mem_counter[4407] = 4'b0000;
    GSharePlugin_logic_mem_counter[4408] = 4'b0000;
    GSharePlugin_logic_mem_counter[4409] = 4'b0000;
    GSharePlugin_logic_mem_counter[4410] = 4'b0000;
    GSharePlugin_logic_mem_counter[4411] = 4'b0000;
    GSharePlugin_logic_mem_counter[4412] = 4'b0000;
    GSharePlugin_logic_mem_counter[4413] = 4'b0000;
    GSharePlugin_logic_mem_counter[4414] = 4'b0000;
    GSharePlugin_logic_mem_counter[4415] = 4'b0000;
    GSharePlugin_logic_mem_counter[4416] = 4'b0000;
    GSharePlugin_logic_mem_counter[4417] = 4'b0000;
    GSharePlugin_logic_mem_counter[4418] = 4'b0000;
    GSharePlugin_logic_mem_counter[4419] = 4'b0000;
    GSharePlugin_logic_mem_counter[4420] = 4'b0000;
    GSharePlugin_logic_mem_counter[4421] = 4'b0000;
    GSharePlugin_logic_mem_counter[4422] = 4'b0000;
    GSharePlugin_logic_mem_counter[4423] = 4'b0000;
    GSharePlugin_logic_mem_counter[4424] = 4'b0000;
    GSharePlugin_logic_mem_counter[4425] = 4'b0000;
    GSharePlugin_logic_mem_counter[4426] = 4'b0000;
    GSharePlugin_logic_mem_counter[4427] = 4'b0000;
    GSharePlugin_logic_mem_counter[4428] = 4'b0000;
    GSharePlugin_logic_mem_counter[4429] = 4'b0000;
    GSharePlugin_logic_mem_counter[4430] = 4'b0000;
    GSharePlugin_logic_mem_counter[4431] = 4'b0000;
    GSharePlugin_logic_mem_counter[4432] = 4'b0000;
    GSharePlugin_logic_mem_counter[4433] = 4'b0000;
    GSharePlugin_logic_mem_counter[4434] = 4'b0000;
    GSharePlugin_logic_mem_counter[4435] = 4'b0000;
    GSharePlugin_logic_mem_counter[4436] = 4'b0000;
    GSharePlugin_logic_mem_counter[4437] = 4'b0000;
    GSharePlugin_logic_mem_counter[4438] = 4'b0000;
    GSharePlugin_logic_mem_counter[4439] = 4'b0000;
    GSharePlugin_logic_mem_counter[4440] = 4'b0000;
    GSharePlugin_logic_mem_counter[4441] = 4'b0000;
    GSharePlugin_logic_mem_counter[4442] = 4'b0000;
    GSharePlugin_logic_mem_counter[4443] = 4'b0000;
    GSharePlugin_logic_mem_counter[4444] = 4'b0000;
    GSharePlugin_logic_mem_counter[4445] = 4'b0000;
    GSharePlugin_logic_mem_counter[4446] = 4'b0000;
    GSharePlugin_logic_mem_counter[4447] = 4'b0000;
    GSharePlugin_logic_mem_counter[4448] = 4'b0000;
    GSharePlugin_logic_mem_counter[4449] = 4'b0000;
    GSharePlugin_logic_mem_counter[4450] = 4'b0000;
    GSharePlugin_logic_mem_counter[4451] = 4'b0000;
    GSharePlugin_logic_mem_counter[4452] = 4'b0000;
    GSharePlugin_logic_mem_counter[4453] = 4'b0000;
    GSharePlugin_logic_mem_counter[4454] = 4'b0000;
    GSharePlugin_logic_mem_counter[4455] = 4'b0000;
    GSharePlugin_logic_mem_counter[4456] = 4'b0000;
    GSharePlugin_logic_mem_counter[4457] = 4'b0000;
    GSharePlugin_logic_mem_counter[4458] = 4'b0000;
    GSharePlugin_logic_mem_counter[4459] = 4'b0000;
    GSharePlugin_logic_mem_counter[4460] = 4'b0000;
    GSharePlugin_logic_mem_counter[4461] = 4'b0000;
    GSharePlugin_logic_mem_counter[4462] = 4'b0000;
    GSharePlugin_logic_mem_counter[4463] = 4'b0000;
    GSharePlugin_logic_mem_counter[4464] = 4'b0000;
    GSharePlugin_logic_mem_counter[4465] = 4'b0000;
    GSharePlugin_logic_mem_counter[4466] = 4'b0000;
    GSharePlugin_logic_mem_counter[4467] = 4'b0000;
    GSharePlugin_logic_mem_counter[4468] = 4'b0000;
    GSharePlugin_logic_mem_counter[4469] = 4'b0000;
    GSharePlugin_logic_mem_counter[4470] = 4'b0000;
    GSharePlugin_logic_mem_counter[4471] = 4'b0000;
    GSharePlugin_logic_mem_counter[4472] = 4'b0000;
    GSharePlugin_logic_mem_counter[4473] = 4'b0000;
    GSharePlugin_logic_mem_counter[4474] = 4'b0000;
    GSharePlugin_logic_mem_counter[4475] = 4'b0000;
    GSharePlugin_logic_mem_counter[4476] = 4'b0000;
    GSharePlugin_logic_mem_counter[4477] = 4'b0000;
    GSharePlugin_logic_mem_counter[4478] = 4'b0000;
    GSharePlugin_logic_mem_counter[4479] = 4'b0000;
    GSharePlugin_logic_mem_counter[4480] = 4'b0000;
    GSharePlugin_logic_mem_counter[4481] = 4'b0000;
    GSharePlugin_logic_mem_counter[4482] = 4'b0000;
    GSharePlugin_logic_mem_counter[4483] = 4'b0000;
    GSharePlugin_logic_mem_counter[4484] = 4'b0000;
    GSharePlugin_logic_mem_counter[4485] = 4'b0000;
    GSharePlugin_logic_mem_counter[4486] = 4'b0000;
    GSharePlugin_logic_mem_counter[4487] = 4'b0000;
    GSharePlugin_logic_mem_counter[4488] = 4'b0000;
    GSharePlugin_logic_mem_counter[4489] = 4'b0000;
    GSharePlugin_logic_mem_counter[4490] = 4'b0000;
    GSharePlugin_logic_mem_counter[4491] = 4'b0000;
    GSharePlugin_logic_mem_counter[4492] = 4'b0000;
    GSharePlugin_logic_mem_counter[4493] = 4'b0000;
    GSharePlugin_logic_mem_counter[4494] = 4'b0000;
    GSharePlugin_logic_mem_counter[4495] = 4'b0000;
    GSharePlugin_logic_mem_counter[4496] = 4'b0000;
    GSharePlugin_logic_mem_counter[4497] = 4'b0000;
    GSharePlugin_logic_mem_counter[4498] = 4'b0000;
    GSharePlugin_logic_mem_counter[4499] = 4'b0000;
    GSharePlugin_logic_mem_counter[4500] = 4'b0000;
    GSharePlugin_logic_mem_counter[4501] = 4'b0000;
    GSharePlugin_logic_mem_counter[4502] = 4'b0000;
    GSharePlugin_logic_mem_counter[4503] = 4'b0000;
    GSharePlugin_logic_mem_counter[4504] = 4'b0000;
    GSharePlugin_logic_mem_counter[4505] = 4'b0000;
    GSharePlugin_logic_mem_counter[4506] = 4'b0000;
    GSharePlugin_logic_mem_counter[4507] = 4'b0000;
    GSharePlugin_logic_mem_counter[4508] = 4'b0000;
    GSharePlugin_logic_mem_counter[4509] = 4'b0000;
    GSharePlugin_logic_mem_counter[4510] = 4'b0000;
    GSharePlugin_logic_mem_counter[4511] = 4'b0000;
    GSharePlugin_logic_mem_counter[4512] = 4'b0000;
    GSharePlugin_logic_mem_counter[4513] = 4'b0000;
    GSharePlugin_logic_mem_counter[4514] = 4'b0000;
    GSharePlugin_logic_mem_counter[4515] = 4'b0000;
    GSharePlugin_logic_mem_counter[4516] = 4'b0000;
    GSharePlugin_logic_mem_counter[4517] = 4'b0000;
    GSharePlugin_logic_mem_counter[4518] = 4'b0000;
    GSharePlugin_logic_mem_counter[4519] = 4'b0000;
    GSharePlugin_logic_mem_counter[4520] = 4'b0000;
    GSharePlugin_logic_mem_counter[4521] = 4'b0000;
    GSharePlugin_logic_mem_counter[4522] = 4'b0000;
    GSharePlugin_logic_mem_counter[4523] = 4'b0000;
    GSharePlugin_logic_mem_counter[4524] = 4'b0000;
    GSharePlugin_logic_mem_counter[4525] = 4'b0000;
    GSharePlugin_logic_mem_counter[4526] = 4'b0000;
    GSharePlugin_logic_mem_counter[4527] = 4'b0000;
    GSharePlugin_logic_mem_counter[4528] = 4'b0000;
    GSharePlugin_logic_mem_counter[4529] = 4'b0000;
    GSharePlugin_logic_mem_counter[4530] = 4'b0000;
    GSharePlugin_logic_mem_counter[4531] = 4'b0000;
    GSharePlugin_logic_mem_counter[4532] = 4'b0000;
    GSharePlugin_logic_mem_counter[4533] = 4'b0000;
    GSharePlugin_logic_mem_counter[4534] = 4'b0000;
    GSharePlugin_logic_mem_counter[4535] = 4'b0000;
    GSharePlugin_logic_mem_counter[4536] = 4'b0000;
    GSharePlugin_logic_mem_counter[4537] = 4'b0000;
    GSharePlugin_logic_mem_counter[4538] = 4'b0000;
    GSharePlugin_logic_mem_counter[4539] = 4'b0000;
    GSharePlugin_logic_mem_counter[4540] = 4'b0000;
    GSharePlugin_logic_mem_counter[4541] = 4'b0000;
    GSharePlugin_logic_mem_counter[4542] = 4'b0000;
    GSharePlugin_logic_mem_counter[4543] = 4'b0000;
    GSharePlugin_logic_mem_counter[4544] = 4'b0000;
    GSharePlugin_logic_mem_counter[4545] = 4'b0000;
    GSharePlugin_logic_mem_counter[4546] = 4'b0000;
    GSharePlugin_logic_mem_counter[4547] = 4'b0000;
    GSharePlugin_logic_mem_counter[4548] = 4'b0000;
    GSharePlugin_logic_mem_counter[4549] = 4'b0000;
    GSharePlugin_logic_mem_counter[4550] = 4'b0000;
    GSharePlugin_logic_mem_counter[4551] = 4'b0000;
    GSharePlugin_logic_mem_counter[4552] = 4'b0000;
    GSharePlugin_logic_mem_counter[4553] = 4'b0000;
    GSharePlugin_logic_mem_counter[4554] = 4'b0000;
    GSharePlugin_logic_mem_counter[4555] = 4'b0000;
    GSharePlugin_logic_mem_counter[4556] = 4'b0000;
    GSharePlugin_logic_mem_counter[4557] = 4'b0000;
    GSharePlugin_logic_mem_counter[4558] = 4'b0000;
    GSharePlugin_logic_mem_counter[4559] = 4'b0000;
    GSharePlugin_logic_mem_counter[4560] = 4'b0000;
    GSharePlugin_logic_mem_counter[4561] = 4'b0000;
    GSharePlugin_logic_mem_counter[4562] = 4'b0000;
    GSharePlugin_logic_mem_counter[4563] = 4'b0000;
    GSharePlugin_logic_mem_counter[4564] = 4'b0000;
    GSharePlugin_logic_mem_counter[4565] = 4'b0000;
    GSharePlugin_logic_mem_counter[4566] = 4'b0000;
    GSharePlugin_logic_mem_counter[4567] = 4'b0000;
    GSharePlugin_logic_mem_counter[4568] = 4'b0000;
    GSharePlugin_logic_mem_counter[4569] = 4'b0000;
    GSharePlugin_logic_mem_counter[4570] = 4'b0000;
    GSharePlugin_logic_mem_counter[4571] = 4'b0000;
    GSharePlugin_logic_mem_counter[4572] = 4'b0000;
    GSharePlugin_logic_mem_counter[4573] = 4'b0000;
    GSharePlugin_logic_mem_counter[4574] = 4'b0000;
    GSharePlugin_logic_mem_counter[4575] = 4'b0000;
    GSharePlugin_logic_mem_counter[4576] = 4'b0000;
    GSharePlugin_logic_mem_counter[4577] = 4'b0000;
    GSharePlugin_logic_mem_counter[4578] = 4'b0000;
    GSharePlugin_logic_mem_counter[4579] = 4'b0000;
    GSharePlugin_logic_mem_counter[4580] = 4'b0000;
    GSharePlugin_logic_mem_counter[4581] = 4'b0000;
    GSharePlugin_logic_mem_counter[4582] = 4'b0000;
    GSharePlugin_logic_mem_counter[4583] = 4'b0000;
    GSharePlugin_logic_mem_counter[4584] = 4'b0000;
    GSharePlugin_logic_mem_counter[4585] = 4'b0000;
    GSharePlugin_logic_mem_counter[4586] = 4'b0000;
    GSharePlugin_logic_mem_counter[4587] = 4'b0000;
    GSharePlugin_logic_mem_counter[4588] = 4'b0000;
    GSharePlugin_logic_mem_counter[4589] = 4'b0000;
    GSharePlugin_logic_mem_counter[4590] = 4'b0000;
    GSharePlugin_logic_mem_counter[4591] = 4'b0000;
    GSharePlugin_logic_mem_counter[4592] = 4'b0000;
    GSharePlugin_logic_mem_counter[4593] = 4'b0000;
    GSharePlugin_logic_mem_counter[4594] = 4'b0000;
    GSharePlugin_logic_mem_counter[4595] = 4'b0000;
    GSharePlugin_logic_mem_counter[4596] = 4'b0000;
    GSharePlugin_logic_mem_counter[4597] = 4'b0000;
    GSharePlugin_logic_mem_counter[4598] = 4'b0000;
    GSharePlugin_logic_mem_counter[4599] = 4'b0000;
    GSharePlugin_logic_mem_counter[4600] = 4'b0000;
    GSharePlugin_logic_mem_counter[4601] = 4'b0000;
    GSharePlugin_logic_mem_counter[4602] = 4'b0000;
    GSharePlugin_logic_mem_counter[4603] = 4'b0000;
    GSharePlugin_logic_mem_counter[4604] = 4'b0000;
    GSharePlugin_logic_mem_counter[4605] = 4'b0000;
    GSharePlugin_logic_mem_counter[4606] = 4'b0000;
    GSharePlugin_logic_mem_counter[4607] = 4'b0000;
    GSharePlugin_logic_mem_counter[4608] = 4'b0000;
    GSharePlugin_logic_mem_counter[4609] = 4'b0000;
    GSharePlugin_logic_mem_counter[4610] = 4'b0000;
    GSharePlugin_logic_mem_counter[4611] = 4'b0000;
    GSharePlugin_logic_mem_counter[4612] = 4'b0000;
    GSharePlugin_logic_mem_counter[4613] = 4'b0000;
    GSharePlugin_logic_mem_counter[4614] = 4'b0000;
    GSharePlugin_logic_mem_counter[4615] = 4'b0000;
    GSharePlugin_logic_mem_counter[4616] = 4'b0000;
    GSharePlugin_logic_mem_counter[4617] = 4'b0000;
    GSharePlugin_logic_mem_counter[4618] = 4'b0000;
    GSharePlugin_logic_mem_counter[4619] = 4'b0000;
    GSharePlugin_logic_mem_counter[4620] = 4'b0000;
    GSharePlugin_logic_mem_counter[4621] = 4'b0000;
    GSharePlugin_logic_mem_counter[4622] = 4'b0000;
    GSharePlugin_logic_mem_counter[4623] = 4'b0000;
    GSharePlugin_logic_mem_counter[4624] = 4'b0000;
    GSharePlugin_logic_mem_counter[4625] = 4'b0000;
    GSharePlugin_logic_mem_counter[4626] = 4'b0000;
    GSharePlugin_logic_mem_counter[4627] = 4'b0000;
    GSharePlugin_logic_mem_counter[4628] = 4'b0000;
    GSharePlugin_logic_mem_counter[4629] = 4'b0000;
    GSharePlugin_logic_mem_counter[4630] = 4'b0000;
    GSharePlugin_logic_mem_counter[4631] = 4'b0000;
    GSharePlugin_logic_mem_counter[4632] = 4'b0000;
    GSharePlugin_logic_mem_counter[4633] = 4'b0000;
    GSharePlugin_logic_mem_counter[4634] = 4'b0000;
    GSharePlugin_logic_mem_counter[4635] = 4'b0000;
    GSharePlugin_logic_mem_counter[4636] = 4'b0000;
    GSharePlugin_logic_mem_counter[4637] = 4'b0000;
    GSharePlugin_logic_mem_counter[4638] = 4'b0000;
    GSharePlugin_logic_mem_counter[4639] = 4'b0000;
    GSharePlugin_logic_mem_counter[4640] = 4'b0000;
    GSharePlugin_logic_mem_counter[4641] = 4'b0000;
    GSharePlugin_logic_mem_counter[4642] = 4'b0000;
    GSharePlugin_logic_mem_counter[4643] = 4'b0000;
    GSharePlugin_logic_mem_counter[4644] = 4'b0000;
    GSharePlugin_logic_mem_counter[4645] = 4'b0000;
    GSharePlugin_logic_mem_counter[4646] = 4'b0000;
    GSharePlugin_logic_mem_counter[4647] = 4'b0000;
    GSharePlugin_logic_mem_counter[4648] = 4'b0000;
    GSharePlugin_logic_mem_counter[4649] = 4'b0000;
    GSharePlugin_logic_mem_counter[4650] = 4'b0000;
    GSharePlugin_logic_mem_counter[4651] = 4'b0000;
    GSharePlugin_logic_mem_counter[4652] = 4'b0000;
    GSharePlugin_logic_mem_counter[4653] = 4'b0000;
    GSharePlugin_logic_mem_counter[4654] = 4'b0000;
    GSharePlugin_logic_mem_counter[4655] = 4'b0000;
    GSharePlugin_logic_mem_counter[4656] = 4'b0000;
    GSharePlugin_logic_mem_counter[4657] = 4'b0000;
    GSharePlugin_logic_mem_counter[4658] = 4'b0000;
    GSharePlugin_logic_mem_counter[4659] = 4'b0000;
    GSharePlugin_logic_mem_counter[4660] = 4'b0000;
    GSharePlugin_logic_mem_counter[4661] = 4'b0000;
    GSharePlugin_logic_mem_counter[4662] = 4'b0000;
    GSharePlugin_logic_mem_counter[4663] = 4'b0000;
    GSharePlugin_logic_mem_counter[4664] = 4'b0000;
    GSharePlugin_logic_mem_counter[4665] = 4'b0000;
    GSharePlugin_logic_mem_counter[4666] = 4'b0000;
    GSharePlugin_logic_mem_counter[4667] = 4'b0000;
    GSharePlugin_logic_mem_counter[4668] = 4'b0000;
    GSharePlugin_logic_mem_counter[4669] = 4'b0000;
    GSharePlugin_logic_mem_counter[4670] = 4'b0000;
    GSharePlugin_logic_mem_counter[4671] = 4'b0000;
    GSharePlugin_logic_mem_counter[4672] = 4'b0000;
    GSharePlugin_logic_mem_counter[4673] = 4'b0000;
    GSharePlugin_logic_mem_counter[4674] = 4'b0000;
    GSharePlugin_logic_mem_counter[4675] = 4'b0000;
    GSharePlugin_logic_mem_counter[4676] = 4'b0000;
    GSharePlugin_logic_mem_counter[4677] = 4'b0000;
    GSharePlugin_logic_mem_counter[4678] = 4'b0000;
    GSharePlugin_logic_mem_counter[4679] = 4'b0000;
    GSharePlugin_logic_mem_counter[4680] = 4'b0000;
    GSharePlugin_logic_mem_counter[4681] = 4'b0000;
    GSharePlugin_logic_mem_counter[4682] = 4'b0000;
    GSharePlugin_logic_mem_counter[4683] = 4'b0000;
    GSharePlugin_logic_mem_counter[4684] = 4'b0000;
    GSharePlugin_logic_mem_counter[4685] = 4'b0000;
    GSharePlugin_logic_mem_counter[4686] = 4'b0000;
    GSharePlugin_logic_mem_counter[4687] = 4'b0000;
    GSharePlugin_logic_mem_counter[4688] = 4'b0000;
    GSharePlugin_logic_mem_counter[4689] = 4'b0000;
    GSharePlugin_logic_mem_counter[4690] = 4'b0000;
    GSharePlugin_logic_mem_counter[4691] = 4'b0000;
    GSharePlugin_logic_mem_counter[4692] = 4'b0000;
    GSharePlugin_logic_mem_counter[4693] = 4'b0000;
    GSharePlugin_logic_mem_counter[4694] = 4'b0000;
    GSharePlugin_logic_mem_counter[4695] = 4'b0000;
    GSharePlugin_logic_mem_counter[4696] = 4'b0000;
    GSharePlugin_logic_mem_counter[4697] = 4'b0000;
    GSharePlugin_logic_mem_counter[4698] = 4'b0000;
    GSharePlugin_logic_mem_counter[4699] = 4'b0000;
    GSharePlugin_logic_mem_counter[4700] = 4'b0000;
    GSharePlugin_logic_mem_counter[4701] = 4'b0000;
    GSharePlugin_logic_mem_counter[4702] = 4'b0000;
    GSharePlugin_logic_mem_counter[4703] = 4'b0000;
    GSharePlugin_logic_mem_counter[4704] = 4'b0000;
    GSharePlugin_logic_mem_counter[4705] = 4'b0000;
    GSharePlugin_logic_mem_counter[4706] = 4'b0000;
    GSharePlugin_logic_mem_counter[4707] = 4'b0000;
    GSharePlugin_logic_mem_counter[4708] = 4'b0000;
    GSharePlugin_logic_mem_counter[4709] = 4'b0000;
    GSharePlugin_logic_mem_counter[4710] = 4'b0000;
    GSharePlugin_logic_mem_counter[4711] = 4'b0000;
    GSharePlugin_logic_mem_counter[4712] = 4'b0000;
    GSharePlugin_logic_mem_counter[4713] = 4'b0000;
    GSharePlugin_logic_mem_counter[4714] = 4'b0000;
    GSharePlugin_logic_mem_counter[4715] = 4'b0000;
    GSharePlugin_logic_mem_counter[4716] = 4'b0000;
    GSharePlugin_logic_mem_counter[4717] = 4'b0000;
    GSharePlugin_logic_mem_counter[4718] = 4'b0000;
    GSharePlugin_logic_mem_counter[4719] = 4'b0000;
    GSharePlugin_logic_mem_counter[4720] = 4'b0000;
    GSharePlugin_logic_mem_counter[4721] = 4'b0000;
    GSharePlugin_logic_mem_counter[4722] = 4'b0000;
    GSharePlugin_logic_mem_counter[4723] = 4'b0000;
    GSharePlugin_logic_mem_counter[4724] = 4'b0000;
    GSharePlugin_logic_mem_counter[4725] = 4'b0000;
    GSharePlugin_logic_mem_counter[4726] = 4'b0000;
    GSharePlugin_logic_mem_counter[4727] = 4'b0000;
    GSharePlugin_logic_mem_counter[4728] = 4'b0000;
    GSharePlugin_logic_mem_counter[4729] = 4'b0000;
    GSharePlugin_logic_mem_counter[4730] = 4'b0000;
    GSharePlugin_logic_mem_counter[4731] = 4'b0000;
    GSharePlugin_logic_mem_counter[4732] = 4'b0000;
    GSharePlugin_logic_mem_counter[4733] = 4'b0000;
    GSharePlugin_logic_mem_counter[4734] = 4'b0000;
    GSharePlugin_logic_mem_counter[4735] = 4'b0000;
    GSharePlugin_logic_mem_counter[4736] = 4'b0000;
    GSharePlugin_logic_mem_counter[4737] = 4'b0000;
    GSharePlugin_logic_mem_counter[4738] = 4'b0000;
    GSharePlugin_logic_mem_counter[4739] = 4'b0000;
    GSharePlugin_logic_mem_counter[4740] = 4'b0000;
    GSharePlugin_logic_mem_counter[4741] = 4'b0000;
    GSharePlugin_logic_mem_counter[4742] = 4'b0000;
    GSharePlugin_logic_mem_counter[4743] = 4'b0000;
    GSharePlugin_logic_mem_counter[4744] = 4'b0000;
    GSharePlugin_logic_mem_counter[4745] = 4'b0000;
    GSharePlugin_logic_mem_counter[4746] = 4'b0000;
    GSharePlugin_logic_mem_counter[4747] = 4'b0000;
    GSharePlugin_logic_mem_counter[4748] = 4'b0000;
    GSharePlugin_logic_mem_counter[4749] = 4'b0000;
    GSharePlugin_logic_mem_counter[4750] = 4'b0000;
    GSharePlugin_logic_mem_counter[4751] = 4'b0000;
    GSharePlugin_logic_mem_counter[4752] = 4'b0000;
    GSharePlugin_logic_mem_counter[4753] = 4'b0000;
    GSharePlugin_logic_mem_counter[4754] = 4'b0000;
    GSharePlugin_logic_mem_counter[4755] = 4'b0000;
    GSharePlugin_logic_mem_counter[4756] = 4'b0000;
    GSharePlugin_logic_mem_counter[4757] = 4'b0000;
    GSharePlugin_logic_mem_counter[4758] = 4'b0000;
    GSharePlugin_logic_mem_counter[4759] = 4'b0000;
    GSharePlugin_logic_mem_counter[4760] = 4'b0000;
    GSharePlugin_logic_mem_counter[4761] = 4'b0000;
    GSharePlugin_logic_mem_counter[4762] = 4'b0000;
    GSharePlugin_logic_mem_counter[4763] = 4'b0000;
    GSharePlugin_logic_mem_counter[4764] = 4'b0000;
    GSharePlugin_logic_mem_counter[4765] = 4'b0000;
    GSharePlugin_logic_mem_counter[4766] = 4'b0000;
    GSharePlugin_logic_mem_counter[4767] = 4'b0000;
    GSharePlugin_logic_mem_counter[4768] = 4'b0000;
    GSharePlugin_logic_mem_counter[4769] = 4'b0000;
    GSharePlugin_logic_mem_counter[4770] = 4'b0000;
    GSharePlugin_logic_mem_counter[4771] = 4'b0000;
    GSharePlugin_logic_mem_counter[4772] = 4'b0000;
    GSharePlugin_logic_mem_counter[4773] = 4'b0000;
    GSharePlugin_logic_mem_counter[4774] = 4'b0000;
    GSharePlugin_logic_mem_counter[4775] = 4'b0000;
    GSharePlugin_logic_mem_counter[4776] = 4'b0000;
    GSharePlugin_logic_mem_counter[4777] = 4'b0000;
    GSharePlugin_logic_mem_counter[4778] = 4'b0000;
    GSharePlugin_logic_mem_counter[4779] = 4'b0000;
    GSharePlugin_logic_mem_counter[4780] = 4'b0000;
    GSharePlugin_logic_mem_counter[4781] = 4'b0000;
    GSharePlugin_logic_mem_counter[4782] = 4'b0000;
    GSharePlugin_logic_mem_counter[4783] = 4'b0000;
    GSharePlugin_logic_mem_counter[4784] = 4'b0000;
    GSharePlugin_logic_mem_counter[4785] = 4'b0000;
    GSharePlugin_logic_mem_counter[4786] = 4'b0000;
    GSharePlugin_logic_mem_counter[4787] = 4'b0000;
    GSharePlugin_logic_mem_counter[4788] = 4'b0000;
    GSharePlugin_logic_mem_counter[4789] = 4'b0000;
    GSharePlugin_logic_mem_counter[4790] = 4'b0000;
    GSharePlugin_logic_mem_counter[4791] = 4'b0000;
    GSharePlugin_logic_mem_counter[4792] = 4'b0000;
    GSharePlugin_logic_mem_counter[4793] = 4'b0000;
    GSharePlugin_logic_mem_counter[4794] = 4'b0000;
    GSharePlugin_logic_mem_counter[4795] = 4'b0000;
    GSharePlugin_logic_mem_counter[4796] = 4'b0000;
    GSharePlugin_logic_mem_counter[4797] = 4'b0000;
    GSharePlugin_logic_mem_counter[4798] = 4'b0000;
    GSharePlugin_logic_mem_counter[4799] = 4'b0000;
    GSharePlugin_logic_mem_counter[4800] = 4'b0000;
    GSharePlugin_logic_mem_counter[4801] = 4'b0000;
    GSharePlugin_logic_mem_counter[4802] = 4'b0000;
    GSharePlugin_logic_mem_counter[4803] = 4'b0000;
    GSharePlugin_logic_mem_counter[4804] = 4'b0000;
    GSharePlugin_logic_mem_counter[4805] = 4'b0000;
    GSharePlugin_logic_mem_counter[4806] = 4'b0000;
    GSharePlugin_logic_mem_counter[4807] = 4'b0000;
    GSharePlugin_logic_mem_counter[4808] = 4'b0000;
    GSharePlugin_logic_mem_counter[4809] = 4'b0000;
    GSharePlugin_logic_mem_counter[4810] = 4'b0000;
    GSharePlugin_logic_mem_counter[4811] = 4'b0000;
    GSharePlugin_logic_mem_counter[4812] = 4'b0000;
    GSharePlugin_logic_mem_counter[4813] = 4'b0000;
    GSharePlugin_logic_mem_counter[4814] = 4'b0000;
    GSharePlugin_logic_mem_counter[4815] = 4'b0000;
    GSharePlugin_logic_mem_counter[4816] = 4'b0000;
    GSharePlugin_logic_mem_counter[4817] = 4'b0000;
    GSharePlugin_logic_mem_counter[4818] = 4'b0000;
    GSharePlugin_logic_mem_counter[4819] = 4'b0000;
    GSharePlugin_logic_mem_counter[4820] = 4'b0000;
    GSharePlugin_logic_mem_counter[4821] = 4'b0000;
    GSharePlugin_logic_mem_counter[4822] = 4'b0000;
    GSharePlugin_logic_mem_counter[4823] = 4'b0000;
    GSharePlugin_logic_mem_counter[4824] = 4'b0000;
    GSharePlugin_logic_mem_counter[4825] = 4'b0000;
    GSharePlugin_logic_mem_counter[4826] = 4'b0000;
    GSharePlugin_logic_mem_counter[4827] = 4'b0000;
    GSharePlugin_logic_mem_counter[4828] = 4'b0000;
    GSharePlugin_logic_mem_counter[4829] = 4'b0000;
    GSharePlugin_logic_mem_counter[4830] = 4'b0000;
    GSharePlugin_logic_mem_counter[4831] = 4'b0000;
    GSharePlugin_logic_mem_counter[4832] = 4'b0000;
    GSharePlugin_logic_mem_counter[4833] = 4'b0000;
    GSharePlugin_logic_mem_counter[4834] = 4'b0000;
    GSharePlugin_logic_mem_counter[4835] = 4'b0000;
    GSharePlugin_logic_mem_counter[4836] = 4'b0000;
    GSharePlugin_logic_mem_counter[4837] = 4'b0000;
    GSharePlugin_logic_mem_counter[4838] = 4'b0000;
    GSharePlugin_logic_mem_counter[4839] = 4'b0000;
    GSharePlugin_logic_mem_counter[4840] = 4'b0000;
    GSharePlugin_logic_mem_counter[4841] = 4'b0000;
    GSharePlugin_logic_mem_counter[4842] = 4'b0000;
    GSharePlugin_logic_mem_counter[4843] = 4'b0000;
    GSharePlugin_logic_mem_counter[4844] = 4'b0000;
    GSharePlugin_logic_mem_counter[4845] = 4'b0000;
    GSharePlugin_logic_mem_counter[4846] = 4'b0000;
    GSharePlugin_logic_mem_counter[4847] = 4'b0000;
    GSharePlugin_logic_mem_counter[4848] = 4'b0000;
    GSharePlugin_logic_mem_counter[4849] = 4'b0000;
    GSharePlugin_logic_mem_counter[4850] = 4'b0000;
    GSharePlugin_logic_mem_counter[4851] = 4'b0000;
    GSharePlugin_logic_mem_counter[4852] = 4'b0000;
    GSharePlugin_logic_mem_counter[4853] = 4'b0000;
    GSharePlugin_logic_mem_counter[4854] = 4'b0000;
    GSharePlugin_logic_mem_counter[4855] = 4'b0000;
    GSharePlugin_logic_mem_counter[4856] = 4'b0000;
    GSharePlugin_logic_mem_counter[4857] = 4'b0000;
    GSharePlugin_logic_mem_counter[4858] = 4'b0000;
    GSharePlugin_logic_mem_counter[4859] = 4'b0000;
    GSharePlugin_logic_mem_counter[4860] = 4'b0000;
    GSharePlugin_logic_mem_counter[4861] = 4'b0000;
    GSharePlugin_logic_mem_counter[4862] = 4'b0000;
    GSharePlugin_logic_mem_counter[4863] = 4'b0000;
    GSharePlugin_logic_mem_counter[4864] = 4'b0000;
    GSharePlugin_logic_mem_counter[4865] = 4'b0000;
    GSharePlugin_logic_mem_counter[4866] = 4'b0000;
    GSharePlugin_logic_mem_counter[4867] = 4'b0000;
    GSharePlugin_logic_mem_counter[4868] = 4'b0000;
    GSharePlugin_logic_mem_counter[4869] = 4'b0000;
    GSharePlugin_logic_mem_counter[4870] = 4'b0000;
    GSharePlugin_logic_mem_counter[4871] = 4'b0000;
    GSharePlugin_logic_mem_counter[4872] = 4'b0000;
    GSharePlugin_logic_mem_counter[4873] = 4'b0000;
    GSharePlugin_logic_mem_counter[4874] = 4'b0000;
    GSharePlugin_logic_mem_counter[4875] = 4'b0000;
    GSharePlugin_logic_mem_counter[4876] = 4'b0000;
    GSharePlugin_logic_mem_counter[4877] = 4'b0000;
    GSharePlugin_logic_mem_counter[4878] = 4'b0000;
    GSharePlugin_logic_mem_counter[4879] = 4'b0000;
    GSharePlugin_logic_mem_counter[4880] = 4'b0000;
    GSharePlugin_logic_mem_counter[4881] = 4'b0000;
    GSharePlugin_logic_mem_counter[4882] = 4'b0000;
    GSharePlugin_logic_mem_counter[4883] = 4'b0000;
    GSharePlugin_logic_mem_counter[4884] = 4'b0000;
    GSharePlugin_logic_mem_counter[4885] = 4'b0000;
    GSharePlugin_logic_mem_counter[4886] = 4'b0000;
    GSharePlugin_logic_mem_counter[4887] = 4'b0000;
    GSharePlugin_logic_mem_counter[4888] = 4'b0000;
    GSharePlugin_logic_mem_counter[4889] = 4'b0000;
    GSharePlugin_logic_mem_counter[4890] = 4'b0000;
    GSharePlugin_logic_mem_counter[4891] = 4'b0000;
    GSharePlugin_logic_mem_counter[4892] = 4'b0000;
    GSharePlugin_logic_mem_counter[4893] = 4'b0000;
    GSharePlugin_logic_mem_counter[4894] = 4'b0000;
    GSharePlugin_logic_mem_counter[4895] = 4'b0000;
    GSharePlugin_logic_mem_counter[4896] = 4'b0000;
    GSharePlugin_logic_mem_counter[4897] = 4'b0000;
    GSharePlugin_logic_mem_counter[4898] = 4'b0000;
    GSharePlugin_logic_mem_counter[4899] = 4'b0000;
    GSharePlugin_logic_mem_counter[4900] = 4'b0000;
    GSharePlugin_logic_mem_counter[4901] = 4'b0000;
    GSharePlugin_logic_mem_counter[4902] = 4'b0000;
    GSharePlugin_logic_mem_counter[4903] = 4'b0000;
    GSharePlugin_logic_mem_counter[4904] = 4'b0000;
    GSharePlugin_logic_mem_counter[4905] = 4'b0000;
    GSharePlugin_logic_mem_counter[4906] = 4'b0000;
    GSharePlugin_logic_mem_counter[4907] = 4'b0000;
    GSharePlugin_logic_mem_counter[4908] = 4'b0000;
    GSharePlugin_logic_mem_counter[4909] = 4'b0000;
    GSharePlugin_logic_mem_counter[4910] = 4'b0000;
    GSharePlugin_logic_mem_counter[4911] = 4'b0000;
    GSharePlugin_logic_mem_counter[4912] = 4'b0000;
    GSharePlugin_logic_mem_counter[4913] = 4'b0000;
    GSharePlugin_logic_mem_counter[4914] = 4'b0000;
    GSharePlugin_logic_mem_counter[4915] = 4'b0000;
    GSharePlugin_logic_mem_counter[4916] = 4'b0000;
    GSharePlugin_logic_mem_counter[4917] = 4'b0000;
    GSharePlugin_logic_mem_counter[4918] = 4'b0000;
    GSharePlugin_logic_mem_counter[4919] = 4'b0000;
    GSharePlugin_logic_mem_counter[4920] = 4'b0000;
    GSharePlugin_logic_mem_counter[4921] = 4'b0000;
    GSharePlugin_logic_mem_counter[4922] = 4'b0000;
    GSharePlugin_logic_mem_counter[4923] = 4'b0000;
    GSharePlugin_logic_mem_counter[4924] = 4'b0000;
    GSharePlugin_logic_mem_counter[4925] = 4'b0000;
    GSharePlugin_logic_mem_counter[4926] = 4'b0000;
    GSharePlugin_logic_mem_counter[4927] = 4'b0000;
    GSharePlugin_logic_mem_counter[4928] = 4'b0000;
    GSharePlugin_logic_mem_counter[4929] = 4'b0000;
    GSharePlugin_logic_mem_counter[4930] = 4'b0000;
    GSharePlugin_logic_mem_counter[4931] = 4'b0000;
    GSharePlugin_logic_mem_counter[4932] = 4'b0000;
    GSharePlugin_logic_mem_counter[4933] = 4'b0000;
    GSharePlugin_logic_mem_counter[4934] = 4'b0000;
    GSharePlugin_logic_mem_counter[4935] = 4'b0000;
    GSharePlugin_logic_mem_counter[4936] = 4'b0000;
    GSharePlugin_logic_mem_counter[4937] = 4'b0000;
    GSharePlugin_logic_mem_counter[4938] = 4'b0000;
    GSharePlugin_logic_mem_counter[4939] = 4'b0000;
    GSharePlugin_logic_mem_counter[4940] = 4'b0000;
    GSharePlugin_logic_mem_counter[4941] = 4'b0000;
    GSharePlugin_logic_mem_counter[4942] = 4'b0000;
    GSharePlugin_logic_mem_counter[4943] = 4'b0000;
    GSharePlugin_logic_mem_counter[4944] = 4'b0000;
    GSharePlugin_logic_mem_counter[4945] = 4'b0000;
    GSharePlugin_logic_mem_counter[4946] = 4'b0000;
    GSharePlugin_logic_mem_counter[4947] = 4'b0000;
    GSharePlugin_logic_mem_counter[4948] = 4'b0000;
    GSharePlugin_logic_mem_counter[4949] = 4'b0000;
    GSharePlugin_logic_mem_counter[4950] = 4'b0000;
    GSharePlugin_logic_mem_counter[4951] = 4'b0000;
    GSharePlugin_logic_mem_counter[4952] = 4'b0000;
    GSharePlugin_logic_mem_counter[4953] = 4'b0000;
    GSharePlugin_logic_mem_counter[4954] = 4'b0000;
    GSharePlugin_logic_mem_counter[4955] = 4'b0000;
    GSharePlugin_logic_mem_counter[4956] = 4'b0000;
    GSharePlugin_logic_mem_counter[4957] = 4'b0000;
    GSharePlugin_logic_mem_counter[4958] = 4'b0000;
    GSharePlugin_logic_mem_counter[4959] = 4'b0000;
    GSharePlugin_logic_mem_counter[4960] = 4'b0000;
    GSharePlugin_logic_mem_counter[4961] = 4'b0000;
    GSharePlugin_logic_mem_counter[4962] = 4'b0000;
    GSharePlugin_logic_mem_counter[4963] = 4'b0000;
    GSharePlugin_logic_mem_counter[4964] = 4'b0000;
    GSharePlugin_logic_mem_counter[4965] = 4'b0000;
    GSharePlugin_logic_mem_counter[4966] = 4'b0000;
    GSharePlugin_logic_mem_counter[4967] = 4'b0000;
    GSharePlugin_logic_mem_counter[4968] = 4'b0000;
    GSharePlugin_logic_mem_counter[4969] = 4'b0000;
    GSharePlugin_logic_mem_counter[4970] = 4'b0000;
    GSharePlugin_logic_mem_counter[4971] = 4'b0000;
    GSharePlugin_logic_mem_counter[4972] = 4'b0000;
    GSharePlugin_logic_mem_counter[4973] = 4'b0000;
    GSharePlugin_logic_mem_counter[4974] = 4'b0000;
    GSharePlugin_logic_mem_counter[4975] = 4'b0000;
    GSharePlugin_logic_mem_counter[4976] = 4'b0000;
    GSharePlugin_logic_mem_counter[4977] = 4'b0000;
    GSharePlugin_logic_mem_counter[4978] = 4'b0000;
    GSharePlugin_logic_mem_counter[4979] = 4'b0000;
    GSharePlugin_logic_mem_counter[4980] = 4'b0000;
    GSharePlugin_logic_mem_counter[4981] = 4'b0000;
    GSharePlugin_logic_mem_counter[4982] = 4'b0000;
    GSharePlugin_logic_mem_counter[4983] = 4'b0000;
    GSharePlugin_logic_mem_counter[4984] = 4'b0000;
    GSharePlugin_logic_mem_counter[4985] = 4'b0000;
    GSharePlugin_logic_mem_counter[4986] = 4'b0000;
    GSharePlugin_logic_mem_counter[4987] = 4'b0000;
    GSharePlugin_logic_mem_counter[4988] = 4'b0000;
    GSharePlugin_logic_mem_counter[4989] = 4'b0000;
    GSharePlugin_logic_mem_counter[4990] = 4'b0000;
    GSharePlugin_logic_mem_counter[4991] = 4'b0000;
    GSharePlugin_logic_mem_counter[4992] = 4'b0000;
    GSharePlugin_logic_mem_counter[4993] = 4'b0000;
    GSharePlugin_logic_mem_counter[4994] = 4'b0000;
    GSharePlugin_logic_mem_counter[4995] = 4'b0000;
    GSharePlugin_logic_mem_counter[4996] = 4'b0000;
    GSharePlugin_logic_mem_counter[4997] = 4'b0000;
    GSharePlugin_logic_mem_counter[4998] = 4'b0000;
    GSharePlugin_logic_mem_counter[4999] = 4'b0000;
    GSharePlugin_logic_mem_counter[5000] = 4'b0000;
    GSharePlugin_logic_mem_counter[5001] = 4'b0000;
    GSharePlugin_logic_mem_counter[5002] = 4'b0000;
    GSharePlugin_logic_mem_counter[5003] = 4'b0000;
    GSharePlugin_logic_mem_counter[5004] = 4'b0000;
    GSharePlugin_logic_mem_counter[5005] = 4'b0000;
    GSharePlugin_logic_mem_counter[5006] = 4'b0000;
    GSharePlugin_logic_mem_counter[5007] = 4'b0000;
    GSharePlugin_logic_mem_counter[5008] = 4'b0000;
    GSharePlugin_logic_mem_counter[5009] = 4'b0000;
    GSharePlugin_logic_mem_counter[5010] = 4'b0000;
    GSharePlugin_logic_mem_counter[5011] = 4'b0000;
    GSharePlugin_logic_mem_counter[5012] = 4'b0000;
    GSharePlugin_logic_mem_counter[5013] = 4'b0000;
    GSharePlugin_logic_mem_counter[5014] = 4'b0000;
    GSharePlugin_logic_mem_counter[5015] = 4'b0000;
    GSharePlugin_logic_mem_counter[5016] = 4'b0000;
    GSharePlugin_logic_mem_counter[5017] = 4'b0000;
    GSharePlugin_logic_mem_counter[5018] = 4'b0000;
    GSharePlugin_logic_mem_counter[5019] = 4'b0000;
    GSharePlugin_logic_mem_counter[5020] = 4'b0000;
    GSharePlugin_logic_mem_counter[5021] = 4'b0000;
    GSharePlugin_logic_mem_counter[5022] = 4'b0000;
    GSharePlugin_logic_mem_counter[5023] = 4'b0000;
    GSharePlugin_logic_mem_counter[5024] = 4'b0000;
    GSharePlugin_logic_mem_counter[5025] = 4'b0000;
    GSharePlugin_logic_mem_counter[5026] = 4'b0000;
    GSharePlugin_logic_mem_counter[5027] = 4'b0000;
    GSharePlugin_logic_mem_counter[5028] = 4'b0000;
    GSharePlugin_logic_mem_counter[5029] = 4'b0000;
    GSharePlugin_logic_mem_counter[5030] = 4'b0000;
    GSharePlugin_logic_mem_counter[5031] = 4'b0000;
    GSharePlugin_logic_mem_counter[5032] = 4'b0000;
    GSharePlugin_logic_mem_counter[5033] = 4'b0000;
    GSharePlugin_logic_mem_counter[5034] = 4'b0000;
    GSharePlugin_logic_mem_counter[5035] = 4'b0000;
    GSharePlugin_logic_mem_counter[5036] = 4'b0000;
    GSharePlugin_logic_mem_counter[5037] = 4'b0000;
    GSharePlugin_logic_mem_counter[5038] = 4'b0000;
    GSharePlugin_logic_mem_counter[5039] = 4'b0000;
    GSharePlugin_logic_mem_counter[5040] = 4'b0000;
    GSharePlugin_logic_mem_counter[5041] = 4'b0000;
    GSharePlugin_logic_mem_counter[5042] = 4'b0000;
    GSharePlugin_logic_mem_counter[5043] = 4'b0000;
    GSharePlugin_logic_mem_counter[5044] = 4'b0000;
    GSharePlugin_logic_mem_counter[5045] = 4'b0000;
    GSharePlugin_logic_mem_counter[5046] = 4'b0000;
    GSharePlugin_logic_mem_counter[5047] = 4'b0000;
    GSharePlugin_logic_mem_counter[5048] = 4'b0000;
    GSharePlugin_logic_mem_counter[5049] = 4'b0000;
    GSharePlugin_logic_mem_counter[5050] = 4'b0000;
    GSharePlugin_logic_mem_counter[5051] = 4'b0000;
    GSharePlugin_logic_mem_counter[5052] = 4'b0000;
    GSharePlugin_logic_mem_counter[5053] = 4'b0000;
    GSharePlugin_logic_mem_counter[5054] = 4'b0000;
    GSharePlugin_logic_mem_counter[5055] = 4'b0000;
    GSharePlugin_logic_mem_counter[5056] = 4'b0000;
    GSharePlugin_logic_mem_counter[5057] = 4'b0000;
    GSharePlugin_logic_mem_counter[5058] = 4'b0000;
    GSharePlugin_logic_mem_counter[5059] = 4'b0000;
    GSharePlugin_logic_mem_counter[5060] = 4'b0000;
    GSharePlugin_logic_mem_counter[5061] = 4'b0000;
    GSharePlugin_logic_mem_counter[5062] = 4'b0000;
    GSharePlugin_logic_mem_counter[5063] = 4'b0000;
    GSharePlugin_logic_mem_counter[5064] = 4'b0000;
    GSharePlugin_logic_mem_counter[5065] = 4'b0000;
    GSharePlugin_logic_mem_counter[5066] = 4'b0000;
    GSharePlugin_logic_mem_counter[5067] = 4'b0000;
    GSharePlugin_logic_mem_counter[5068] = 4'b0000;
    GSharePlugin_logic_mem_counter[5069] = 4'b0000;
    GSharePlugin_logic_mem_counter[5070] = 4'b0000;
    GSharePlugin_logic_mem_counter[5071] = 4'b0000;
    GSharePlugin_logic_mem_counter[5072] = 4'b0000;
    GSharePlugin_logic_mem_counter[5073] = 4'b0000;
    GSharePlugin_logic_mem_counter[5074] = 4'b0000;
    GSharePlugin_logic_mem_counter[5075] = 4'b0000;
    GSharePlugin_logic_mem_counter[5076] = 4'b0000;
    GSharePlugin_logic_mem_counter[5077] = 4'b0000;
    GSharePlugin_logic_mem_counter[5078] = 4'b0000;
    GSharePlugin_logic_mem_counter[5079] = 4'b0000;
    GSharePlugin_logic_mem_counter[5080] = 4'b0000;
    GSharePlugin_logic_mem_counter[5081] = 4'b0000;
    GSharePlugin_logic_mem_counter[5082] = 4'b0000;
    GSharePlugin_logic_mem_counter[5083] = 4'b0000;
    GSharePlugin_logic_mem_counter[5084] = 4'b0000;
    GSharePlugin_logic_mem_counter[5085] = 4'b0000;
    GSharePlugin_logic_mem_counter[5086] = 4'b0000;
    GSharePlugin_logic_mem_counter[5087] = 4'b0000;
    GSharePlugin_logic_mem_counter[5088] = 4'b0000;
    GSharePlugin_logic_mem_counter[5089] = 4'b0000;
    GSharePlugin_logic_mem_counter[5090] = 4'b0000;
    GSharePlugin_logic_mem_counter[5091] = 4'b0000;
    GSharePlugin_logic_mem_counter[5092] = 4'b0000;
    GSharePlugin_logic_mem_counter[5093] = 4'b0000;
    GSharePlugin_logic_mem_counter[5094] = 4'b0000;
    GSharePlugin_logic_mem_counter[5095] = 4'b0000;
    GSharePlugin_logic_mem_counter[5096] = 4'b0000;
    GSharePlugin_logic_mem_counter[5097] = 4'b0000;
    GSharePlugin_logic_mem_counter[5098] = 4'b0000;
    GSharePlugin_logic_mem_counter[5099] = 4'b0000;
    GSharePlugin_logic_mem_counter[5100] = 4'b0000;
    GSharePlugin_logic_mem_counter[5101] = 4'b0000;
    GSharePlugin_logic_mem_counter[5102] = 4'b0000;
    GSharePlugin_logic_mem_counter[5103] = 4'b0000;
    GSharePlugin_logic_mem_counter[5104] = 4'b0000;
    GSharePlugin_logic_mem_counter[5105] = 4'b0000;
    GSharePlugin_logic_mem_counter[5106] = 4'b0000;
    GSharePlugin_logic_mem_counter[5107] = 4'b0000;
    GSharePlugin_logic_mem_counter[5108] = 4'b0000;
    GSharePlugin_logic_mem_counter[5109] = 4'b0000;
    GSharePlugin_logic_mem_counter[5110] = 4'b0000;
    GSharePlugin_logic_mem_counter[5111] = 4'b0000;
    GSharePlugin_logic_mem_counter[5112] = 4'b0000;
    GSharePlugin_logic_mem_counter[5113] = 4'b0000;
    GSharePlugin_logic_mem_counter[5114] = 4'b0000;
    GSharePlugin_logic_mem_counter[5115] = 4'b0000;
    GSharePlugin_logic_mem_counter[5116] = 4'b0000;
    GSharePlugin_logic_mem_counter[5117] = 4'b0000;
    GSharePlugin_logic_mem_counter[5118] = 4'b0000;
    GSharePlugin_logic_mem_counter[5119] = 4'b0000;
    GSharePlugin_logic_mem_counter[5120] = 4'b0000;
    GSharePlugin_logic_mem_counter[5121] = 4'b0000;
    GSharePlugin_logic_mem_counter[5122] = 4'b0000;
    GSharePlugin_logic_mem_counter[5123] = 4'b0000;
    GSharePlugin_logic_mem_counter[5124] = 4'b0000;
    GSharePlugin_logic_mem_counter[5125] = 4'b0000;
    GSharePlugin_logic_mem_counter[5126] = 4'b0000;
    GSharePlugin_logic_mem_counter[5127] = 4'b0000;
    GSharePlugin_logic_mem_counter[5128] = 4'b0000;
    GSharePlugin_logic_mem_counter[5129] = 4'b0000;
    GSharePlugin_logic_mem_counter[5130] = 4'b0000;
    GSharePlugin_logic_mem_counter[5131] = 4'b0000;
    GSharePlugin_logic_mem_counter[5132] = 4'b0000;
    GSharePlugin_logic_mem_counter[5133] = 4'b0000;
    GSharePlugin_logic_mem_counter[5134] = 4'b0000;
    GSharePlugin_logic_mem_counter[5135] = 4'b0000;
    GSharePlugin_logic_mem_counter[5136] = 4'b0000;
    GSharePlugin_logic_mem_counter[5137] = 4'b0000;
    GSharePlugin_logic_mem_counter[5138] = 4'b0000;
    GSharePlugin_logic_mem_counter[5139] = 4'b0000;
    GSharePlugin_logic_mem_counter[5140] = 4'b0000;
    GSharePlugin_logic_mem_counter[5141] = 4'b0000;
    GSharePlugin_logic_mem_counter[5142] = 4'b0000;
    GSharePlugin_logic_mem_counter[5143] = 4'b0000;
    GSharePlugin_logic_mem_counter[5144] = 4'b0000;
    GSharePlugin_logic_mem_counter[5145] = 4'b0000;
    GSharePlugin_logic_mem_counter[5146] = 4'b0000;
    GSharePlugin_logic_mem_counter[5147] = 4'b0000;
    GSharePlugin_logic_mem_counter[5148] = 4'b0000;
    GSharePlugin_logic_mem_counter[5149] = 4'b0000;
    GSharePlugin_logic_mem_counter[5150] = 4'b0000;
    GSharePlugin_logic_mem_counter[5151] = 4'b0000;
    GSharePlugin_logic_mem_counter[5152] = 4'b0000;
    GSharePlugin_logic_mem_counter[5153] = 4'b0000;
    GSharePlugin_logic_mem_counter[5154] = 4'b0000;
    GSharePlugin_logic_mem_counter[5155] = 4'b0000;
    GSharePlugin_logic_mem_counter[5156] = 4'b0000;
    GSharePlugin_logic_mem_counter[5157] = 4'b0000;
    GSharePlugin_logic_mem_counter[5158] = 4'b0000;
    GSharePlugin_logic_mem_counter[5159] = 4'b0000;
    GSharePlugin_logic_mem_counter[5160] = 4'b0000;
    GSharePlugin_logic_mem_counter[5161] = 4'b0000;
    GSharePlugin_logic_mem_counter[5162] = 4'b0000;
    GSharePlugin_logic_mem_counter[5163] = 4'b0000;
    GSharePlugin_logic_mem_counter[5164] = 4'b0000;
    GSharePlugin_logic_mem_counter[5165] = 4'b0000;
    GSharePlugin_logic_mem_counter[5166] = 4'b0000;
    GSharePlugin_logic_mem_counter[5167] = 4'b0000;
    GSharePlugin_logic_mem_counter[5168] = 4'b0000;
    GSharePlugin_logic_mem_counter[5169] = 4'b0000;
    GSharePlugin_logic_mem_counter[5170] = 4'b0000;
    GSharePlugin_logic_mem_counter[5171] = 4'b0000;
    GSharePlugin_logic_mem_counter[5172] = 4'b0000;
    GSharePlugin_logic_mem_counter[5173] = 4'b0000;
    GSharePlugin_logic_mem_counter[5174] = 4'b0000;
    GSharePlugin_logic_mem_counter[5175] = 4'b0000;
    GSharePlugin_logic_mem_counter[5176] = 4'b0000;
    GSharePlugin_logic_mem_counter[5177] = 4'b0000;
    GSharePlugin_logic_mem_counter[5178] = 4'b0000;
    GSharePlugin_logic_mem_counter[5179] = 4'b0000;
    GSharePlugin_logic_mem_counter[5180] = 4'b0000;
    GSharePlugin_logic_mem_counter[5181] = 4'b0000;
    GSharePlugin_logic_mem_counter[5182] = 4'b0000;
    GSharePlugin_logic_mem_counter[5183] = 4'b0000;
    GSharePlugin_logic_mem_counter[5184] = 4'b0000;
    GSharePlugin_logic_mem_counter[5185] = 4'b0000;
    GSharePlugin_logic_mem_counter[5186] = 4'b0000;
    GSharePlugin_logic_mem_counter[5187] = 4'b0000;
    GSharePlugin_logic_mem_counter[5188] = 4'b0000;
    GSharePlugin_logic_mem_counter[5189] = 4'b0000;
    GSharePlugin_logic_mem_counter[5190] = 4'b0000;
    GSharePlugin_logic_mem_counter[5191] = 4'b0000;
    GSharePlugin_logic_mem_counter[5192] = 4'b0000;
    GSharePlugin_logic_mem_counter[5193] = 4'b0000;
    GSharePlugin_logic_mem_counter[5194] = 4'b0000;
    GSharePlugin_logic_mem_counter[5195] = 4'b0000;
    GSharePlugin_logic_mem_counter[5196] = 4'b0000;
    GSharePlugin_logic_mem_counter[5197] = 4'b0000;
    GSharePlugin_logic_mem_counter[5198] = 4'b0000;
    GSharePlugin_logic_mem_counter[5199] = 4'b0000;
    GSharePlugin_logic_mem_counter[5200] = 4'b0000;
    GSharePlugin_logic_mem_counter[5201] = 4'b0000;
    GSharePlugin_logic_mem_counter[5202] = 4'b0000;
    GSharePlugin_logic_mem_counter[5203] = 4'b0000;
    GSharePlugin_logic_mem_counter[5204] = 4'b0000;
    GSharePlugin_logic_mem_counter[5205] = 4'b0000;
    GSharePlugin_logic_mem_counter[5206] = 4'b0000;
    GSharePlugin_logic_mem_counter[5207] = 4'b0000;
    GSharePlugin_logic_mem_counter[5208] = 4'b0000;
    GSharePlugin_logic_mem_counter[5209] = 4'b0000;
    GSharePlugin_logic_mem_counter[5210] = 4'b0000;
    GSharePlugin_logic_mem_counter[5211] = 4'b0000;
    GSharePlugin_logic_mem_counter[5212] = 4'b0000;
    GSharePlugin_logic_mem_counter[5213] = 4'b0000;
    GSharePlugin_logic_mem_counter[5214] = 4'b0000;
    GSharePlugin_logic_mem_counter[5215] = 4'b0000;
    GSharePlugin_logic_mem_counter[5216] = 4'b0000;
    GSharePlugin_logic_mem_counter[5217] = 4'b0000;
    GSharePlugin_logic_mem_counter[5218] = 4'b0000;
    GSharePlugin_logic_mem_counter[5219] = 4'b0000;
    GSharePlugin_logic_mem_counter[5220] = 4'b0000;
    GSharePlugin_logic_mem_counter[5221] = 4'b0000;
    GSharePlugin_logic_mem_counter[5222] = 4'b0000;
    GSharePlugin_logic_mem_counter[5223] = 4'b0000;
    GSharePlugin_logic_mem_counter[5224] = 4'b0000;
    GSharePlugin_logic_mem_counter[5225] = 4'b0000;
    GSharePlugin_logic_mem_counter[5226] = 4'b0000;
    GSharePlugin_logic_mem_counter[5227] = 4'b0000;
    GSharePlugin_logic_mem_counter[5228] = 4'b0000;
    GSharePlugin_logic_mem_counter[5229] = 4'b0000;
    GSharePlugin_logic_mem_counter[5230] = 4'b0000;
    GSharePlugin_logic_mem_counter[5231] = 4'b0000;
    GSharePlugin_logic_mem_counter[5232] = 4'b0000;
    GSharePlugin_logic_mem_counter[5233] = 4'b0000;
    GSharePlugin_logic_mem_counter[5234] = 4'b0000;
    GSharePlugin_logic_mem_counter[5235] = 4'b0000;
    GSharePlugin_logic_mem_counter[5236] = 4'b0000;
    GSharePlugin_logic_mem_counter[5237] = 4'b0000;
    GSharePlugin_logic_mem_counter[5238] = 4'b0000;
    GSharePlugin_logic_mem_counter[5239] = 4'b0000;
    GSharePlugin_logic_mem_counter[5240] = 4'b0000;
    GSharePlugin_logic_mem_counter[5241] = 4'b0000;
    GSharePlugin_logic_mem_counter[5242] = 4'b0000;
    GSharePlugin_logic_mem_counter[5243] = 4'b0000;
    GSharePlugin_logic_mem_counter[5244] = 4'b0000;
    GSharePlugin_logic_mem_counter[5245] = 4'b0000;
    GSharePlugin_logic_mem_counter[5246] = 4'b0000;
    GSharePlugin_logic_mem_counter[5247] = 4'b0000;
    GSharePlugin_logic_mem_counter[5248] = 4'b0000;
    GSharePlugin_logic_mem_counter[5249] = 4'b0000;
    GSharePlugin_logic_mem_counter[5250] = 4'b0000;
    GSharePlugin_logic_mem_counter[5251] = 4'b0000;
    GSharePlugin_logic_mem_counter[5252] = 4'b0000;
    GSharePlugin_logic_mem_counter[5253] = 4'b0000;
    GSharePlugin_logic_mem_counter[5254] = 4'b0000;
    GSharePlugin_logic_mem_counter[5255] = 4'b0000;
    GSharePlugin_logic_mem_counter[5256] = 4'b0000;
    GSharePlugin_logic_mem_counter[5257] = 4'b0000;
    GSharePlugin_logic_mem_counter[5258] = 4'b0000;
    GSharePlugin_logic_mem_counter[5259] = 4'b0000;
    GSharePlugin_logic_mem_counter[5260] = 4'b0000;
    GSharePlugin_logic_mem_counter[5261] = 4'b0000;
    GSharePlugin_logic_mem_counter[5262] = 4'b0000;
    GSharePlugin_logic_mem_counter[5263] = 4'b0000;
    GSharePlugin_logic_mem_counter[5264] = 4'b0000;
    GSharePlugin_logic_mem_counter[5265] = 4'b0000;
    GSharePlugin_logic_mem_counter[5266] = 4'b0000;
    GSharePlugin_logic_mem_counter[5267] = 4'b0000;
    GSharePlugin_logic_mem_counter[5268] = 4'b0000;
    GSharePlugin_logic_mem_counter[5269] = 4'b0000;
    GSharePlugin_logic_mem_counter[5270] = 4'b0000;
    GSharePlugin_logic_mem_counter[5271] = 4'b0000;
    GSharePlugin_logic_mem_counter[5272] = 4'b0000;
    GSharePlugin_logic_mem_counter[5273] = 4'b0000;
    GSharePlugin_logic_mem_counter[5274] = 4'b0000;
    GSharePlugin_logic_mem_counter[5275] = 4'b0000;
    GSharePlugin_logic_mem_counter[5276] = 4'b0000;
    GSharePlugin_logic_mem_counter[5277] = 4'b0000;
    GSharePlugin_logic_mem_counter[5278] = 4'b0000;
    GSharePlugin_logic_mem_counter[5279] = 4'b0000;
    GSharePlugin_logic_mem_counter[5280] = 4'b0000;
    GSharePlugin_logic_mem_counter[5281] = 4'b0000;
    GSharePlugin_logic_mem_counter[5282] = 4'b0000;
    GSharePlugin_logic_mem_counter[5283] = 4'b0000;
    GSharePlugin_logic_mem_counter[5284] = 4'b0000;
    GSharePlugin_logic_mem_counter[5285] = 4'b0000;
    GSharePlugin_logic_mem_counter[5286] = 4'b0000;
    GSharePlugin_logic_mem_counter[5287] = 4'b0000;
    GSharePlugin_logic_mem_counter[5288] = 4'b0000;
    GSharePlugin_logic_mem_counter[5289] = 4'b0000;
    GSharePlugin_logic_mem_counter[5290] = 4'b0000;
    GSharePlugin_logic_mem_counter[5291] = 4'b0000;
    GSharePlugin_logic_mem_counter[5292] = 4'b0000;
    GSharePlugin_logic_mem_counter[5293] = 4'b0000;
    GSharePlugin_logic_mem_counter[5294] = 4'b0000;
    GSharePlugin_logic_mem_counter[5295] = 4'b0000;
    GSharePlugin_logic_mem_counter[5296] = 4'b0000;
    GSharePlugin_logic_mem_counter[5297] = 4'b0000;
    GSharePlugin_logic_mem_counter[5298] = 4'b0000;
    GSharePlugin_logic_mem_counter[5299] = 4'b0000;
    GSharePlugin_logic_mem_counter[5300] = 4'b0000;
    GSharePlugin_logic_mem_counter[5301] = 4'b0000;
    GSharePlugin_logic_mem_counter[5302] = 4'b0000;
    GSharePlugin_logic_mem_counter[5303] = 4'b0000;
    GSharePlugin_logic_mem_counter[5304] = 4'b0000;
    GSharePlugin_logic_mem_counter[5305] = 4'b0000;
    GSharePlugin_logic_mem_counter[5306] = 4'b0000;
    GSharePlugin_logic_mem_counter[5307] = 4'b0000;
    GSharePlugin_logic_mem_counter[5308] = 4'b0000;
    GSharePlugin_logic_mem_counter[5309] = 4'b0000;
    GSharePlugin_logic_mem_counter[5310] = 4'b0000;
    GSharePlugin_logic_mem_counter[5311] = 4'b0000;
    GSharePlugin_logic_mem_counter[5312] = 4'b0000;
    GSharePlugin_logic_mem_counter[5313] = 4'b0000;
    GSharePlugin_logic_mem_counter[5314] = 4'b0000;
    GSharePlugin_logic_mem_counter[5315] = 4'b0000;
    GSharePlugin_logic_mem_counter[5316] = 4'b0000;
    GSharePlugin_logic_mem_counter[5317] = 4'b0000;
    GSharePlugin_logic_mem_counter[5318] = 4'b0000;
    GSharePlugin_logic_mem_counter[5319] = 4'b0000;
    GSharePlugin_logic_mem_counter[5320] = 4'b0000;
    GSharePlugin_logic_mem_counter[5321] = 4'b0000;
    GSharePlugin_logic_mem_counter[5322] = 4'b0000;
    GSharePlugin_logic_mem_counter[5323] = 4'b0000;
    GSharePlugin_logic_mem_counter[5324] = 4'b0000;
    GSharePlugin_logic_mem_counter[5325] = 4'b0000;
    GSharePlugin_logic_mem_counter[5326] = 4'b0000;
    GSharePlugin_logic_mem_counter[5327] = 4'b0000;
    GSharePlugin_logic_mem_counter[5328] = 4'b0000;
    GSharePlugin_logic_mem_counter[5329] = 4'b0000;
    GSharePlugin_logic_mem_counter[5330] = 4'b0000;
    GSharePlugin_logic_mem_counter[5331] = 4'b0000;
    GSharePlugin_logic_mem_counter[5332] = 4'b0000;
    GSharePlugin_logic_mem_counter[5333] = 4'b0000;
    GSharePlugin_logic_mem_counter[5334] = 4'b0000;
    GSharePlugin_logic_mem_counter[5335] = 4'b0000;
    GSharePlugin_logic_mem_counter[5336] = 4'b0000;
    GSharePlugin_logic_mem_counter[5337] = 4'b0000;
    GSharePlugin_logic_mem_counter[5338] = 4'b0000;
    GSharePlugin_logic_mem_counter[5339] = 4'b0000;
    GSharePlugin_logic_mem_counter[5340] = 4'b0000;
    GSharePlugin_logic_mem_counter[5341] = 4'b0000;
    GSharePlugin_logic_mem_counter[5342] = 4'b0000;
    GSharePlugin_logic_mem_counter[5343] = 4'b0000;
    GSharePlugin_logic_mem_counter[5344] = 4'b0000;
    GSharePlugin_logic_mem_counter[5345] = 4'b0000;
    GSharePlugin_logic_mem_counter[5346] = 4'b0000;
    GSharePlugin_logic_mem_counter[5347] = 4'b0000;
    GSharePlugin_logic_mem_counter[5348] = 4'b0000;
    GSharePlugin_logic_mem_counter[5349] = 4'b0000;
    GSharePlugin_logic_mem_counter[5350] = 4'b0000;
    GSharePlugin_logic_mem_counter[5351] = 4'b0000;
    GSharePlugin_logic_mem_counter[5352] = 4'b0000;
    GSharePlugin_logic_mem_counter[5353] = 4'b0000;
    GSharePlugin_logic_mem_counter[5354] = 4'b0000;
    GSharePlugin_logic_mem_counter[5355] = 4'b0000;
    GSharePlugin_logic_mem_counter[5356] = 4'b0000;
    GSharePlugin_logic_mem_counter[5357] = 4'b0000;
    GSharePlugin_logic_mem_counter[5358] = 4'b0000;
    GSharePlugin_logic_mem_counter[5359] = 4'b0000;
    GSharePlugin_logic_mem_counter[5360] = 4'b0000;
    GSharePlugin_logic_mem_counter[5361] = 4'b0000;
    GSharePlugin_logic_mem_counter[5362] = 4'b0000;
    GSharePlugin_logic_mem_counter[5363] = 4'b0000;
    GSharePlugin_logic_mem_counter[5364] = 4'b0000;
    GSharePlugin_logic_mem_counter[5365] = 4'b0000;
    GSharePlugin_logic_mem_counter[5366] = 4'b0000;
    GSharePlugin_logic_mem_counter[5367] = 4'b0000;
    GSharePlugin_logic_mem_counter[5368] = 4'b0000;
    GSharePlugin_logic_mem_counter[5369] = 4'b0000;
    GSharePlugin_logic_mem_counter[5370] = 4'b0000;
    GSharePlugin_logic_mem_counter[5371] = 4'b0000;
    GSharePlugin_logic_mem_counter[5372] = 4'b0000;
    GSharePlugin_logic_mem_counter[5373] = 4'b0000;
    GSharePlugin_logic_mem_counter[5374] = 4'b0000;
    GSharePlugin_logic_mem_counter[5375] = 4'b0000;
    GSharePlugin_logic_mem_counter[5376] = 4'b0000;
    GSharePlugin_logic_mem_counter[5377] = 4'b0000;
    GSharePlugin_logic_mem_counter[5378] = 4'b0000;
    GSharePlugin_logic_mem_counter[5379] = 4'b0000;
    GSharePlugin_logic_mem_counter[5380] = 4'b0000;
    GSharePlugin_logic_mem_counter[5381] = 4'b0000;
    GSharePlugin_logic_mem_counter[5382] = 4'b0000;
    GSharePlugin_logic_mem_counter[5383] = 4'b0000;
    GSharePlugin_logic_mem_counter[5384] = 4'b0000;
    GSharePlugin_logic_mem_counter[5385] = 4'b0000;
    GSharePlugin_logic_mem_counter[5386] = 4'b0000;
    GSharePlugin_logic_mem_counter[5387] = 4'b0000;
    GSharePlugin_logic_mem_counter[5388] = 4'b0000;
    GSharePlugin_logic_mem_counter[5389] = 4'b0000;
    GSharePlugin_logic_mem_counter[5390] = 4'b0000;
    GSharePlugin_logic_mem_counter[5391] = 4'b0000;
    GSharePlugin_logic_mem_counter[5392] = 4'b0000;
    GSharePlugin_logic_mem_counter[5393] = 4'b0000;
    GSharePlugin_logic_mem_counter[5394] = 4'b0000;
    GSharePlugin_logic_mem_counter[5395] = 4'b0000;
    GSharePlugin_logic_mem_counter[5396] = 4'b0000;
    GSharePlugin_logic_mem_counter[5397] = 4'b0000;
    GSharePlugin_logic_mem_counter[5398] = 4'b0000;
    GSharePlugin_logic_mem_counter[5399] = 4'b0000;
    GSharePlugin_logic_mem_counter[5400] = 4'b0000;
    GSharePlugin_logic_mem_counter[5401] = 4'b0000;
    GSharePlugin_logic_mem_counter[5402] = 4'b0000;
    GSharePlugin_logic_mem_counter[5403] = 4'b0000;
    GSharePlugin_logic_mem_counter[5404] = 4'b0000;
    GSharePlugin_logic_mem_counter[5405] = 4'b0000;
    GSharePlugin_logic_mem_counter[5406] = 4'b0000;
    GSharePlugin_logic_mem_counter[5407] = 4'b0000;
    GSharePlugin_logic_mem_counter[5408] = 4'b0000;
    GSharePlugin_logic_mem_counter[5409] = 4'b0000;
    GSharePlugin_logic_mem_counter[5410] = 4'b0000;
    GSharePlugin_logic_mem_counter[5411] = 4'b0000;
    GSharePlugin_logic_mem_counter[5412] = 4'b0000;
    GSharePlugin_logic_mem_counter[5413] = 4'b0000;
    GSharePlugin_logic_mem_counter[5414] = 4'b0000;
    GSharePlugin_logic_mem_counter[5415] = 4'b0000;
    GSharePlugin_logic_mem_counter[5416] = 4'b0000;
    GSharePlugin_logic_mem_counter[5417] = 4'b0000;
    GSharePlugin_logic_mem_counter[5418] = 4'b0000;
    GSharePlugin_logic_mem_counter[5419] = 4'b0000;
    GSharePlugin_logic_mem_counter[5420] = 4'b0000;
    GSharePlugin_logic_mem_counter[5421] = 4'b0000;
    GSharePlugin_logic_mem_counter[5422] = 4'b0000;
    GSharePlugin_logic_mem_counter[5423] = 4'b0000;
    GSharePlugin_logic_mem_counter[5424] = 4'b0000;
    GSharePlugin_logic_mem_counter[5425] = 4'b0000;
    GSharePlugin_logic_mem_counter[5426] = 4'b0000;
    GSharePlugin_logic_mem_counter[5427] = 4'b0000;
    GSharePlugin_logic_mem_counter[5428] = 4'b0000;
    GSharePlugin_logic_mem_counter[5429] = 4'b0000;
    GSharePlugin_logic_mem_counter[5430] = 4'b0000;
    GSharePlugin_logic_mem_counter[5431] = 4'b0000;
    GSharePlugin_logic_mem_counter[5432] = 4'b0000;
    GSharePlugin_logic_mem_counter[5433] = 4'b0000;
    GSharePlugin_logic_mem_counter[5434] = 4'b0000;
    GSharePlugin_logic_mem_counter[5435] = 4'b0000;
    GSharePlugin_logic_mem_counter[5436] = 4'b0000;
    GSharePlugin_logic_mem_counter[5437] = 4'b0000;
    GSharePlugin_logic_mem_counter[5438] = 4'b0000;
    GSharePlugin_logic_mem_counter[5439] = 4'b0000;
    GSharePlugin_logic_mem_counter[5440] = 4'b0000;
    GSharePlugin_logic_mem_counter[5441] = 4'b0000;
    GSharePlugin_logic_mem_counter[5442] = 4'b0000;
    GSharePlugin_logic_mem_counter[5443] = 4'b0000;
    GSharePlugin_logic_mem_counter[5444] = 4'b0000;
    GSharePlugin_logic_mem_counter[5445] = 4'b0000;
    GSharePlugin_logic_mem_counter[5446] = 4'b0000;
    GSharePlugin_logic_mem_counter[5447] = 4'b0000;
    GSharePlugin_logic_mem_counter[5448] = 4'b0000;
    GSharePlugin_logic_mem_counter[5449] = 4'b0000;
    GSharePlugin_logic_mem_counter[5450] = 4'b0000;
    GSharePlugin_logic_mem_counter[5451] = 4'b0000;
    GSharePlugin_logic_mem_counter[5452] = 4'b0000;
    GSharePlugin_logic_mem_counter[5453] = 4'b0000;
    GSharePlugin_logic_mem_counter[5454] = 4'b0000;
    GSharePlugin_logic_mem_counter[5455] = 4'b0000;
    GSharePlugin_logic_mem_counter[5456] = 4'b0000;
    GSharePlugin_logic_mem_counter[5457] = 4'b0000;
    GSharePlugin_logic_mem_counter[5458] = 4'b0000;
    GSharePlugin_logic_mem_counter[5459] = 4'b0000;
    GSharePlugin_logic_mem_counter[5460] = 4'b0000;
    GSharePlugin_logic_mem_counter[5461] = 4'b0000;
    GSharePlugin_logic_mem_counter[5462] = 4'b0000;
    GSharePlugin_logic_mem_counter[5463] = 4'b0000;
    GSharePlugin_logic_mem_counter[5464] = 4'b0000;
    GSharePlugin_logic_mem_counter[5465] = 4'b0000;
    GSharePlugin_logic_mem_counter[5466] = 4'b0000;
    GSharePlugin_logic_mem_counter[5467] = 4'b0000;
    GSharePlugin_logic_mem_counter[5468] = 4'b0000;
    GSharePlugin_logic_mem_counter[5469] = 4'b0000;
    GSharePlugin_logic_mem_counter[5470] = 4'b0000;
    GSharePlugin_logic_mem_counter[5471] = 4'b0000;
    GSharePlugin_logic_mem_counter[5472] = 4'b0000;
    GSharePlugin_logic_mem_counter[5473] = 4'b0000;
    GSharePlugin_logic_mem_counter[5474] = 4'b0000;
    GSharePlugin_logic_mem_counter[5475] = 4'b0000;
    GSharePlugin_logic_mem_counter[5476] = 4'b0000;
    GSharePlugin_logic_mem_counter[5477] = 4'b0000;
    GSharePlugin_logic_mem_counter[5478] = 4'b0000;
    GSharePlugin_logic_mem_counter[5479] = 4'b0000;
    GSharePlugin_logic_mem_counter[5480] = 4'b0000;
    GSharePlugin_logic_mem_counter[5481] = 4'b0000;
    GSharePlugin_logic_mem_counter[5482] = 4'b0000;
    GSharePlugin_logic_mem_counter[5483] = 4'b0000;
    GSharePlugin_logic_mem_counter[5484] = 4'b0000;
    GSharePlugin_logic_mem_counter[5485] = 4'b0000;
    GSharePlugin_logic_mem_counter[5486] = 4'b0000;
    GSharePlugin_logic_mem_counter[5487] = 4'b0000;
    GSharePlugin_logic_mem_counter[5488] = 4'b0000;
    GSharePlugin_logic_mem_counter[5489] = 4'b0000;
    GSharePlugin_logic_mem_counter[5490] = 4'b0000;
    GSharePlugin_logic_mem_counter[5491] = 4'b0000;
    GSharePlugin_logic_mem_counter[5492] = 4'b0000;
    GSharePlugin_logic_mem_counter[5493] = 4'b0000;
    GSharePlugin_logic_mem_counter[5494] = 4'b0000;
    GSharePlugin_logic_mem_counter[5495] = 4'b0000;
    GSharePlugin_logic_mem_counter[5496] = 4'b0000;
    GSharePlugin_logic_mem_counter[5497] = 4'b0000;
    GSharePlugin_logic_mem_counter[5498] = 4'b0000;
    GSharePlugin_logic_mem_counter[5499] = 4'b0000;
    GSharePlugin_logic_mem_counter[5500] = 4'b0000;
    GSharePlugin_logic_mem_counter[5501] = 4'b0000;
    GSharePlugin_logic_mem_counter[5502] = 4'b0000;
    GSharePlugin_logic_mem_counter[5503] = 4'b0000;
    GSharePlugin_logic_mem_counter[5504] = 4'b0000;
    GSharePlugin_logic_mem_counter[5505] = 4'b0000;
    GSharePlugin_logic_mem_counter[5506] = 4'b0000;
    GSharePlugin_logic_mem_counter[5507] = 4'b0000;
    GSharePlugin_logic_mem_counter[5508] = 4'b0000;
    GSharePlugin_logic_mem_counter[5509] = 4'b0000;
    GSharePlugin_logic_mem_counter[5510] = 4'b0000;
    GSharePlugin_logic_mem_counter[5511] = 4'b0000;
    GSharePlugin_logic_mem_counter[5512] = 4'b0000;
    GSharePlugin_logic_mem_counter[5513] = 4'b0000;
    GSharePlugin_logic_mem_counter[5514] = 4'b0000;
    GSharePlugin_logic_mem_counter[5515] = 4'b0000;
    GSharePlugin_logic_mem_counter[5516] = 4'b0000;
    GSharePlugin_logic_mem_counter[5517] = 4'b0000;
    GSharePlugin_logic_mem_counter[5518] = 4'b0000;
    GSharePlugin_logic_mem_counter[5519] = 4'b0000;
    GSharePlugin_logic_mem_counter[5520] = 4'b0000;
    GSharePlugin_logic_mem_counter[5521] = 4'b0000;
    GSharePlugin_logic_mem_counter[5522] = 4'b0000;
    GSharePlugin_logic_mem_counter[5523] = 4'b0000;
    GSharePlugin_logic_mem_counter[5524] = 4'b0000;
    GSharePlugin_logic_mem_counter[5525] = 4'b0000;
    GSharePlugin_logic_mem_counter[5526] = 4'b0000;
    GSharePlugin_logic_mem_counter[5527] = 4'b0000;
    GSharePlugin_logic_mem_counter[5528] = 4'b0000;
    GSharePlugin_logic_mem_counter[5529] = 4'b0000;
    GSharePlugin_logic_mem_counter[5530] = 4'b0000;
    GSharePlugin_logic_mem_counter[5531] = 4'b0000;
    GSharePlugin_logic_mem_counter[5532] = 4'b0000;
    GSharePlugin_logic_mem_counter[5533] = 4'b0000;
    GSharePlugin_logic_mem_counter[5534] = 4'b0000;
    GSharePlugin_logic_mem_counter[5535] = 4'b0000;
    GSharePlugin_logic_mem_counter[5536] = 4'b0000;
    GSharePlugin_logic_mem_counter[5537] = 4'b0000;
    GSharePlugin_logic_mem_counter[5538] = 4'b0000;
    GSharePlugin_logic_mem_counter[5539] = 4'b0000;
    GSharePlugin_logic_mem_counter[5540] = 4'b0000;
    GSharePlugin_logic_mem_counter[5541] = 4'b0000;
    GSharePlugin_logic_mem_counter[5542] = 4'b0000;
    GSharePlugin_logic_mem_counter[5543] = 4'b0000;
    GSharePlugin_logic_mem_counter[5544] = 4'b0000;
    GSharePlugin_logic_mem_counter[5545] = 4'b0000;
    GSharePlugin_logic_mem_counter[5546] = 4'b0000;
    GSharePlugin_logic_mem_counter[5547] = 4'b0000;
    GSharePlugin_logic_mem_counter[5548] = 4'b0000;
    GSharePlugin_logic_mem_counter[5549] = 4'b0000;
    GSharePlugin_logic_mem_counter[5550] = 4'b0000;
    GSharePlugin_logic_mem_counter[5551] = 4'b0000;
    GSharePlugin_logic_mem_counter[5552] = 4'b0000;
    GSharePlugin_logic_mem_counter[5553] = 4'b0000;
    GSharePlugin_logic_mem_counter[5554] = 4'b0000;
    GSharePlugin_logic_mem_counter[5555] = 4'b0000;
    GSharePlugin_logic_mem_counter[5556] = 4'b0000;
    GSharePlugin_logic_mem_counter[5557] = 4'b0000;
    GSharePlugin_logic_mem_counter[5558] = 4'b0000;
    GSharePlugin_logic_mem_counter[5559] = 4'b0000;
    GSharePlugin_logic_mem_counter[5560] = 4'b0000;
    GSharePlugin_logic_mem_counter[5561] = 4'b0000;
    GSharePlugin_logic_mem_counter[5562] = 4'b0000;
    GSharePlugin_logic_mem_counter[5563] = 4'b0000;
    GSharePlugin_logic_mem_counter[5564] = 4'b0000;
    GSharePlugin_logic_mem_counter[5565] = 4'b0000;
    GSharePlugin_logic_mem_counter[5566] = 4'b0000;
    GSharePlugin_logic_mem_counter[5567] = 4'b0000;
    GSharePlugin_logic_mem_counter[5568] = 4'b0000;
    GSharePlugin_logic_mem_counter[5569] = 4'b0000;
    GSharePlugin_logic_mem_counter[5570] = 4'b0000;
    GSharePlugin_logic_mem_counter[5571] = 4'b0000;
    GSharePlugin_logic_mem_counter[5572] = 4'b0000;
    GSharePlugin_logic_mem_counter[5573] = 4'b0000;
    GSharePlugin_logic_mem_counter[5574] = 4'b0000;
    GSharePlugin_logic_mem_counter[5575] = 4'b0000;
    GSharePlugin_logic_mem_counter[5576] = 4'b0000;
    GSharePlugin_logic_mem_counter[5577] = 4'b0000;
    GSharePlugin_logic_mem_counter[5578] = 4'b0000;
    GSharePlugin_logic_mem_counter[5579] = 4'b0000;
    GSharePlugin_logic_mem_counter[5580] = 4'b0000;
    GSharePlugin_logic_mem_counter[5581] = 4'b0000;
    GSharePlugin_logic_mem_counter[5582] = 4'b0000;
    GSharePlugin_logic_mem_counter[5583] = 4'b0000;
    GSharePlugin_logic_mem_counter[5584] = 4'b0000;
    GSharePlugin_logic_mem_counter[5585] = 4'b0000;
    GSharePlugin_logic_mem_counter[5586] = 4'b0000;
    GSharePlugin_logic_mem_counter[5587] = 4'b0000;
    GSharePlugin_logic_mem_counter[5588] = 4'b0000;
    GSharePlugin_logic_mem_counter[5589] = 4'b0000;
    GSharePlugin_logic_mem_counter[5590] = 4'b0000;
    GSharePlugin_logic_mem_counter[5591] = 4'b0000;
    GSharePlugin_logic_mem_counter[5592] = 4'b0000;
    GSharePlugin_logic_mem_counter[5593] = 4'b0000;
    GSharePlugin_logic_mem_counter[5594] = 4'b0000;
    GSharePlugin_logic_mem_counter[5595] = 4'b0000;
    GSharePlugin_logic_mem_counter[5596] = 4'b0000;
    GSharePlugin_logic_mem_counter[5597] = 4'b0000;
    GSharePlugin_logic_mem_counter[5598] = 4'b0000;
    GSharePlugin_logic_mem_counter[5599] = 4'b0000;
    GSharePlugin_logic_mem_counter[5600] = 4'b0000;
    GSharePlugin_logic_mem_counter[5601] = 4'b0000;
    GSharePlugin_logic_mem_counter[5602] = 4'b0000;
    GSharePlugin_logic_mem_counter[5603] = 4'b0000;
    GSharePlugin_logic_mem_counter[5604] = 4'b0000;
    GSharePlugin_logic_mem_counter[5605] = 4'b0000;
    GSharePlugin_logic_mem_counter[5606] = 4'b0000;
    GSharePlugin_logic_mem_counter[5607] = 4'b0000;
    GSharePlugin_logic_mem_counter[5608] = 4'b0000;
    GSharePlugin_logic_mem_counter[5609] = 4'b0000;
    GSharePlugin_logic_mem_counter[5610] = 4'b0000;
    GSharePlugin_logic_mem_counter[5611] = 4'b0000;
    GSharePlugin_logic_mem_counter[5612] = 4'b0000;
    GSharePlugin_logic_mem_counter[5613] = 4'b0000;
    GSharePlugin_logic_mem_counter[5614] = 4'b0000;
    GSharePlugin_logic_mem_counter[5615] = 4'b0000;
    GSharePlugin_logic_mem_counter[5616] = 4'b0000;
    GSharePlugin_logic_mem_counter[5617] = 4'b0000;
    GSharePlugin_logic_mem_counter[5618] = 4'b0000;
    GSharePlugin_logic_mem_counter[5619] = 4'b0000;
    GSharePlugin_logic_mem_counter[5620] = 4'b0000;
    GSharePlugin_logic_mem_counter[5621] = 4'b0000;
    GSharePlugin_logic_mem_counter[5622] = 4'b0000;
    GSharePlugin_logic_mem_counter[5623] = 4'b0000;
    GSharePlugin_logic_mem_counter[5624] = 4'b0000;
    GSharePlugin_logic_mem_counter[5625] = 4'b0000;
    GSharePlugin_logic_mem_counter[5626] = 4'b0000;
    GSharePlugin_logic_mem_counter[5627] = 4'b0000;
    GSharePlugin_logic_mem_counter[5628] = 4'b0000;
    GSharePlugin_logic_mem_counter[5629] = 4'b0000;
    GSharePlugin_logic_mem_counter[5630] = 4'b0000;
    GSharePlugin_logic_mem_counter[5631] = 4'b0000;
    GSharePlugin_logic_mem_counter[5632] = 4'b0000;
    GSharePlugin_logic_mem_counter[5633] = 4'b0000;
    GSharePlugin_logic_mem_counter[5634] = 4'b0000;
    GSharePlugin_logic_mem_counter[5635] = 4'b0000;
    GSharePlugin_logic_mem_counter[5636] = 4'b0000;
    GSharePlugin_logic_mem_counter[5637] = 4'b0000;
    GSharePlugin_logic_mem_counter[5638] = 4'b0000;
    GSharePlugin_logic_mem_counter[5639] = 4'b0000;
    GSharePlugin_logic_mem_counter[5640] = 4'b0000;
    GSharePlugin_logic_mem_counter[5641] = 4'b0000;
    GSharePlugin_logic_mem_counter[5642] = 4'b0000;
    GSharePlugin_logic_mem_counter[5643] = 4'b0000;
    GSharePlugin_logic_mem_counter[5644] = 4'b0000;
    GSharePlugin_logic_mem_counter[5645] = 4'b0000;
    GSharePlugin_logic_mem_counter[5646] = 4'b0000;
    GSharePlugin_logic_mem_counter[5647] = 4'b0000;
    GSharePlugin_logic_mem_counter[5648] = 4'b0000;
    GSharePlugin_logic_mem_counter[5649] = 4'b0000;
    GSharePlugin_logic_mem_counter[5650] = 4'b0000;
    GSharePlugin_logic_mem_counter[5651] = 4'b0000;
    GSharePlugin_logic_mem_counter[5652] = 4'b0000;
    GSharePlugin_logic_mem_counter[5653] = 4'b0000;
    GSharePlugin_logic_mem_counter[5654] = 4'b0000;
    GSharePlugin_logic_mem_counter[5655] = 4'b0000;
    GSharePlugin_logic_mem_counter[5656] = 4'b0000;
    GSharePlugin_logic_mem_counter[5657] = 4'b0000;
    GSharePlugin_logic_mem_counter[5658] = 4'b0000;
    GSharePlugin_logic_mem_counter[5659] = 4'b0000;
    GSharePlugin_logic_mem_counter[5660] = 4'b0000;
    GSharePlugin_logic_mem_counter[5661] = 4'b0000;
    GSharePlugin_logic_mem_counter[5662] = 4'b0000;
    GSharePlugin_logic_mem_counter[5663] = 4'b0000;
    GSharePlugin_logic_mem_counter[5664] = 4'b0000;
    GSharePlugin_logic_mem_counter[5665] = 4'b0000;
    GSharePlugin_logic_mem_counter[5666] = 4'b0000;
    GSharePlugin_logic_mem_counter[5667] = 4'b0000;
    GSharePlugin_logic_mem_counter[5668] = 4'b0000;
    GSharePlugin_logic_mem_counter[5669] = 4'b0000;
    GSharePlugin_logic_mem_counter[5670] = 4'b0000;
    GSharePlugin_logic_mem_counter[5671] = 4'b0000;
    GSharePlugin_logic_mem_counter[5672] = 4'b0000;
    GSharePlugin_logic_mem_counter[5673] = 4'b0000;
    GSharePlugin_logic_mem_counter[5674] = 4'b0000;
    GSharePlugin_logic_mem_counter[5675] = 4'b0000;
    GSharePlugin_logic_mem_counter[5676] = 4'b0000;
    GSharePlugin_logic_mem_counter[5677] = 4'b0000;
    GSharePlugin_logic_mem_counter[5678] = 4'b0000;
    GSharePlugin_logic_mem_counter[5679] = 4'b0000;
    GSharePlugin_logic_mem_counter[5680] = 4'b0000;
    GSharePlugin_logic_mem_counter[5681] = 4'b0000;
    GSharePlugin_logic_mem_counter[5682] = 4'b0000;
    GSharePlugin_logic_mem_counter[5683] = 4'b0000;
    GSharePlugin_logic_mem_counter[5684] = 4'b0000;
    GSharePlugin_logic_mem_counter[5685] = 4'b0000;
    GSharePlugin_logic_mem_counter[5686] = 4'b0000;
    GSharePlugin_logic_mem_counter[5687] = 4'b0000;
    GSharePlugin_logic_mem_counter[5688] = 4'b0000;
    GSharePlugin_logic_mem_counter[5689] = 4'b0000;
    GSharePlugin_logic_mem_counter[5690] = 4'b0000;
    GSharePlugin_logic_mem_counter[5691] = 4'b0000;
    GSharePlugin_logic_mem_counter[5692] = 4'b0000;
    GSharePlugin_logic_mem_counter[5693] = 4'b0000;
    GSharePlugin_logic_mem_counter[5694] = 4'b0000;
    GSharePlugin_logic_mem_counter[5695] = 4'b0000;
    GSharePlugin_logic_mem_counter[5696] = 4'b0000;
    GSharePlugin_logic_mem_counter[5697] = 4'b0000;
    GSharePlugin_logic_mem_counter[5698] = 4'b0000;
    GSharePlugin_logic_mem_counter[5699] = 4'b0000;
    GSharePlugin_logic_mem_counter[5700] = 4'b0000;
    GSharePlugin_logic_mem_counter[5701] = 4'b0000;
    GSharePlugin_logic_mem_counter[5702] = 4'b0000;
    GSharePlugin_logic_mem_counter[5703] = 4'b0000;
    GSharePlugin_logic_mem_counter[5704] = 4'b0000;
    GSharePlugin_logic_mem_counter[5705] = 4'b0000;
    GSharePlugin_logic_mem_counter[5706] = 4'b0000;
    GSharePlugin_logic_mem_counter[5707] = 4'b0000;
    GSharePlugin_logic_mem_counter[5708] = 4'b0000;
    GSharePlugin_logic_mem_counter[5709] = 4'b0000;
    GSharePlugin_logic_mem_counter[5710] = 4'b0000;
    GSharePlugin_logic_mem_counter[5711] = 4'b0000;
    GSharePlugin_logic_mem_counter[5712] = 4'b0000;
    GSharePlugin_logic_mem_counter[5713] = 4'b0000;
    GSharePlugin_logic_mem_counter[5714] = 4'b0000;
    GSharePlugin_logic_mem_counter[5715] = 4'b0000;
    GSharePlugin_logic_mem_counter[5716] = 4'b0000;
    GSharePlugin_logic_mem_counter[5717] = 4'b0000;
    GSharePlugin_logic_mem_counter[5718] = 4'b0000;
    GSharePlugin_logic_mem_counter[5719] = 4'b0000;
    GSharePlugin_logic_mem_counter[5720] = 4'b0000;
    GSharePlugin_logic_mem_counter[5721] = 4'b0000;
    GSharePlugin_logic_mem_counter[5722] = 4'b0000;
    GSharePlugin_logic_mem_counter[5723] = 4'b0000;
    GSharePlugin_logic_mem_counter[5724] = 4'b0000;
    GSharePlugin_logic_mem_counter[5725] = 4'b0000;
    GSharePlugin_logic_mem_counter[5726] = 4'b0000;
    GSharePlugin_logic_mem_counter[5727] = 4'b0000;
    GSharePlugin_logic_mem_counter[5728] = 4'b0000;
    GSharePlugin_logic_mem_counter[5729] = 4'b0000;
    GSharePlugin_logic_mem_counter[5730] = 4'b0000;
    GSharePlugin_logic_mem_counter[5731] = 4'b0000;
    GSharePlugin_logic_mem_counter[5732] = 4'b0000;
    GSharePlugin_logic_mem_counter[5733] = 4'b0000;
    GSharePlugin_logic_mem_counter[5734] = 4'b0000;
    GSharePlugin_logic_mem_counter[5735] = 4'b0000;
    GSharePlugin_logic_mem_counter[5736] = 4'b0000;
    GSharePlugin_logic_mem_counter[5737] = 4'b0000;
    GSharePlugin_logic_mem_counter[5738] = 4'b0000;
    GSharePlugin_logic_mem_counter[5739] = 4'b0000;
    GSharePlugin_logic_mem_counter[5740] = 4'b0000;
    GSharePlugin_logic_mem_counter[5741] = 4'b0000;
    GSharePlugin_logic_mem_counter[5742] = 4'b0000;
    GSharePlugin_logic_mem_counter[5743] = 4'b0000;
    GSharePlugin_logic_mem_counter[5744] = 4'b0000;
    GSharePlugin_logic_mem_counter[5745] = 4'b0000;
    GSharePlugin_logic_mem_counter[5746] = 4'b0000;
    GSharePlugin_logic_mem_counter[5747] = 4'b0000;
    GSharePlugin_logic_mem_counter[5748] = 4'b0000;
    GSharePlugin_logic_mem_counter[5749] = 4'b0000;
    GSharePlugin_logic_mem_counter[5750] = 4'b0000;
    GSharePlugin_logic_mem_counter[5751] = 4'b0000;
    GSharePlugin_logic_mem_counter[5752] = 4'b0000;
    GSharePlugin_logic_mem_counter[5753] = 4'b0000;
    GSharePlugin_logic_mem_counter[5754] = 4'b0000;
    GSharePlugin_logic_mem_counter[5755] = 4'b0000;
    GSharePlugin_logic_mem_counter[5756] = 4'b0000;
    GSharePlugin_logic_mem_counter[5757] = 4'b0000;
    GSharePlugin_logic_mem_counter[5758] = 4'b0000;
    GSharePlugin_logic_mem_counter[5759] = 4'b0000;
    GSharePlugin_logic_mem_counter[5760] = 4'b0000;
    GSharePlugin_logic_mem_counter[5761] = 4'b0000;
    GSharePlugin_logic_mem_counter[5762] = 4'b0000;
    GSharePlugin_logic_mem_counter[5763] = 4'b0000;
    GSharePlugin_logic_mem_counter[5764] = 4'b0000;
    GSharePlugin_logic_mem_counter[5765] = 4'b0000;
    GSharePlugin_logic_mem_counter[5766] = 4'b0000;
    GSharePlugin_logic_mem_counter[5767] = 4'b0000;
    GSharePlugin_logic_mem_counter[5768] = 4'b0000;
    GSharePlugin_logic_mem_counter[5769] = 4'b0000;
    GSharePlugin_logic_mem_counter[5770] = 4'b0000;
    GSharePlugin_logic_mem_counter[5771] = 4'b0000;
    GSharePlugin_logic_mem_counter[5772] = 4'b0000;
    GSharePlugin_logic_mem_counter[5773] = 4'b0000;
    GSharePlugin_logic_mem_counter[5774] = 4'b0000;
    GSharePlugin_logic_mem_counter[5775] = 4'b0000;
    GSharePlugin_logic_mem_counter[5776] = 4'b0000;
    GSharePlugin_logic_mem_counter[5777] = 4'b0000;
    GSharePlugin_logic_mem_counter[5778] = 4'b0000;
    GSharePlugin_logic_mem_counter[5779] = 4'b0000;
    GSharePlugin_logic_mem_counter[5780] = 4'b0000;
    GSharePlugin_logic_mem_counter[5781] = 4'b0000;
    GSharePlugin_logic_mem_counter[5782] = 4'b0000;
    GSharePlugin_logic_mem_counter[5783] = 4'b0000;
    GSharePlugin_logic_mem_counter[5784] = 4'b0000;
    GSharePlugin_logic_mem_counter[5785] = 4'b0000;
    GSharePlugin_logic_mem_counter[5786] = 4'b0000;
    GSharePlugin_logic_mem_counter[5787] = 4'b0000;
    GSharePlugin_logic_mem_counter[5788] = 4'b0000;
    GSharePlugin_logic_mem_counter[5789] = 4'b0000;
    GSharePlugin_logic_mem_counter[5790] = 4'b0000;
    GSharePlugin_logic_mem_counter[5791] = 4'b0000;
    GSharePlugin_logic_mem_counter[5792] = 4'b0000;
    GSharePlugin_logic_mem_counter[5793] = 4'b0000;
    GSharePlugin_logic_mem_counter[5794] = 4'b0000;
    GSharePlugin_logic_mem_counter[5795] = 4'b0000;
    GSharePlugin_logic_mem_counter[5796] = 4'b0000;
    GSharePlugin_logic_mem_counter[5797] = 4'b0000;
    GSharePlugin_logic_mem_counter[5798] = 4'b0000;
    GSharePlugin_logic_mem_counter[5799] = 4'b0000;
    GSharePlugin_logic_mem_counter[5800] = 4'b0000;
    GSharePlugin_logic_mem_counter[5801] = 4'b0000;
    GSharePlugin_logic_mem_counter[5802] = 4'b0000;
    GSharePlugin_logic_mem_counter[5803] = 4'b0000;
    GSharePlugin_logic_mem_counter[5804] = 4'b0000;
    GSharePlugin_logic_mem_counter[5805] = 4'b0000;
    GSharePlugin_logic_mem_counter[5806] = 4'b0000;
    GSharePlugin_logic_mem_counter[5807] = 4'b0000;
    GSharePlugin_logic_mem_counter[5808] = 4'b0000;
    GSharePlugin_logic_mem_counter[5809] = 4'b0000;
    GSharePlugin_logic_mem_counter[5810] = 4'b0000;
    GSharePlugin_logic_mem_counter[5811] = 4'b0000;
    GSharePlugin_logic_mem_counter[5812] = 4'b0000;
    GSharePlugin_logic_mem_counter[5813] = 4'b0000;
    GSharePlugin_logic_mem_counter[5814] = 4'b0000;
    GSharePlugin_logic_mem_counter[5815] = 4'b0000;
    GSharePlugin_logic_mem_counter[5816] = 4'b0000;
    GSharePlugin_logic_mem_counter[5817] = 4'b0000;
    GSharePlugin_logic_mem_counter[5818] = 4'b0000;
    GSharePlugin_logic_mem_counter[5819] = 4'b0000;
    GSharePlugin_logic_mem_counter[5820] = 4'b0000;
    GSharePlugin_logic_mem_counter[5821] = 4'b0000;
    GSharePlugin_logic_mem_counter[5822] = 4'b0000;
    GSharePlugin_logic_mem_counter[5823] = 4'b0000;
    GSharePlugin_logic_mem_counter[5824] = 4'b0000;
    GSharePlugin_logic_mem_counter[5825] = 4'b0000;
    GSharePlugin_logic_mem_counter[5826] = 4'b0000;
    GSharePlugin_logic_mem_counter[5827] = 4'b0000;
    GSharePlugin_logic_mem_counter[5828] = 4'b0000;
    GSharePlugin_logic_mem_counter[5829] = 4'b0000;
    GSharePlugin_logic_mem_counter[5830] = 4'b0000;
    GSharePlugin_logic_mem_counter[5831] = 4'b0000;
    GSharePlugin_logic_mem_counter[5832] = 4'b0000;
    GSharePlugin_logic_mem_counter[5833] = 4'b0000;
    GSharePlugin_logic_mem_counter[5834] = 4'b0000;
    GSharePlugin_logic_mem_counter[5835] = 4'b0000;
    GSharePlugin_logic_mem_counter[5836] = 4'b0000;
    GSharePlugin_logic_mem_counter[5837] = 4'b0000;
    GSharePlugin_logic_mem_counter[5838] = 4'b0000;
    GSharePlugin_logic_mem_counter[5839] = 4'b0000;
    GSharePlugin_logic_mem_counter[5840] = 4'b0000;
    GSharePlugin_logic_mem_counter[5841] = 4'b0000;
    GSharePlugin_logic_mem_counter[5842] = 4'b0000;
    GSharePlugin_logic_mem_counter[5843] = 4'b0000;
    GSharePlugin_logic_mem_counter[5844] = 4'b0000;
    GSharePlugin_logic_mem_counter[5845] = 4'b0000;
    GSharePlugin_logic_mem_counter[5846] = 4'b0000;
    GSharePlugin_logic_mem_counter[5847] = 4'b0000;
    GSharePlugin_logic_mem_counter[5848] = 4'b0000;
    GSharePlugin_logic_mem_counter[5849] = 4'b0000;
    GSharePlugin_logic_mem_counter[5850] = 4'b0000;
    GSharePlugin_logic_mem_counter[5851] = 4'b0000;
    GSharePlugin_logic_mem_counter[5852] = 4'b0000;
    GSharePlugin_logic_mem_counter[5853] = 4'b0000;
    GSharePlugin_logic_mem_counter[5854] = 4'b0000;
    GSharePlugin_logic_mem_counter[5855] = 4'b0000;
    GSharePlugin_logic_mem_counter[5856] = 4'b0000;
    GSharePlugin_logic_mem_counter[5857] = 4'b0000;
    GSharePlugin_logic_mem_counter[5858] = 4'b0000;
    GSharePlugin_logic_mem_counter[5859] = 4'b0000;
    GSharePlugin_logic_mem_counter[5860] = 4'b0000;
    GSharePlugin_logic_mem_counter[5861] = 4'b0000;
    GSharePlugin_logic_mem_counter[5862] = 4'b0000;
    GSharePlugin_logic_mem_counter[5863] = 4'b0000;
    GSharePlugin_logic_mem_counter[5864] = 4'b0000;
    GSharePlugin_logic_mem_counter[5865] = 4'b0000;
    GSharePlugin_logic_mem_counter[5866] = 4'b0000;
    GSharePlugin_logic_mem_counter[5867] = 4'b0000;
    GSharePlugin_logic_mem_counter[5868] = 4'b0000;
    GSharePlugin_logic_mem_counter[5869] = 4'b0000;
    GSharePlugin_logic_mem_counter[5870] = 4'b0000;
    GSharePlugin_logic_mem_counter[5871] = 4'b0000;
    GSharePlugin_logic_mem_counter[5872] = 4'b0000;
    GSharePlugin_logic_mem_counter[5873] = 4'b0000;
    GSharePlugin_logic_mem_counter[5874] = 4'b0000;
    GSharePlugin_logic_mem_counter[5875] = 4'b0000;
    GSharePlugin_logic_mem_counter[5876] = 4'b0000;
    GSharePlugin_logic_mem_counter[5877] = 4'b0000;
    GSharePlugin_logic_mem_counter[5878] = 4'b0000;
    GSharePlugin_logic_mem_counter[5879] = 4'b0000;
    GSharePlugin_logic_mem_counter[5880] = 4'b0000;
    GSharePlugin_logic_mem_counter[5881] = 4'b0000;
    GSharePlugin_logic_mem_counter[5882] = 4'b0000;
    GSharePlugin_logic_mem_counter[5883] = 4'b0000;
    GSharePlugin_logic_mem_counter[5884] = 4'b0000;
    GSharePlugin_logic_mem_counter[5885] = 4'b0000;
    GSharePlugin_logic_mem_counter[5886] = 4'b0000;
    GSharePlugin_logic_mem_counter[5887] = 4'b0000;
    GSharePlugin_logic_mem_counter[5888] = 4'b0000;
    GSharePlugin_logic_mem_counter[5889] = 4'b0000;
    GSharePlugin_logic_mem_counter[5890] = 4'b0000;
    GSharePlugin_logic_mem_counter[5891] = 4'b0000;
    GSharePlugin_logic_mem_counter[5892] = 4'b0000;
    GSharePlugin_logic_mem_counter[5893] = 4'b0000;
    GSharePlugin_logic_mem_counter[5894] = 4'b0000;
    GSharePlugin_logic_mem_counter[5895] = 4'b0000;
    GSharePlugin_logic_mem_counter[5896] = 4'b0000;
    GSharePlugin_logic_mem_counter[5897] = 4'b0000;
    GSharePlugin_logic_mem_counter[5898] = 4'b0000;
    GSharePlugin_logic_mem_counter[5899] = 4'b0000;
    GSharePlugin_logic_mem_counter[5900] = 4'b0000;
    GSharePlugin_logic_mem_counter[5901] = 4'b0000;
    GSharePlugin_logic_mem_counter[5902] = 4'b0000;
    GSharePlugin_logic_mem_counter[5903] = 4'b0000;
    GSharePlugin_logic_mem_counter[5904] = 4'b0000;
    GSharePlugin_logic_mem_counter[5905] = 4'b0000;
    GSharePlugin_logic_mem_counter[5906] = 4'b0000;
    GSharePlugin_logic_mem_counter[5907] = 4'b0000;
    GSharePlugin_logic_mem_counter[5908] = 4'b0000;
    GSharePlugin_logic_mem_counter[5909] = 4'b0000;
    GSharePlugin_logic_mem_counter[5910] = 4'b0000;
    GSharePlugin_logic_mem_counter[5911] = 4'b0000;
    GSharePlugin_logic_mem_counter[5912] = 4'b0000;
    GSharePlugin_logic_mem_counter[5913] = 4'b0000;
    GSharePlugin_logic_mem_counter[5914] = 4'b0000;
    GSharePlugin_logic_mem_counter[5915] = 4'b0000;
    GSharePlugin_logic_mem_counter[5916] = 4'b0000;
    GSharePlugin_logic_mem_counter[5917] = 4'b0000;
    GSharePlugin_logic_mem_counter[5918] = 4'b0000;
    GSharePlugin_logic_mem_counter[5919] = 4'b0000;
    GSharePlugin_logic_mem_counter[5920] = 4'b0000;
    GSharePlugin_logic_mem_counter[5921] = 4'b0000;
    GSharePlugin_logic_mem_counter[5922] = 4'b0000;
    GSharePlugin_logic_mem_counter[5923] = 4'b0000;
    GSharePlugin_logic_mem_counter[5924] = 4'b0000;
    GSharePlugin_logic_mem_counter[5925] = 4'b0000;
    GSharePlugin_logic_mem_counter[5926] = 4'b0000;
    GSharePlugin_logic_mem_counter[5927] = 4'b0000;
    GSharePlugin_logic_mem_counter[5928] = 4'b0000;
    GSharePlugin_logic_mem_counter[5929] = 4'b0000;
    GSharePlugin_logic_mem_counter[5930] = 4'b0000;
    GSharePlugin_logic_mem_counter[5931] = 4'b0000;
    GSharePlugin_logic_mem_counter[5932] = 4'b0000;
    GSharePlugin_logic_mem_counter[5933] = 4'b0000;
    GSharePlugin_logic_mem_counter[5934] = 4'b0000;
    GSharePlugin_logic_mem_counter[5935] = 4'b0000;
    GSharePlugin_logic_mem_counter[5936] = 4'b0000;
    GSharePlugin_logic_mem_counter[5937] = 4'b0000;
    GSharePlugin_logic_mem_counter[5938] = 4'b0000;
    GSharePlugin_logic_mem_counter[5939] = 4'b0000;
    GSharePlugin_logic_mem_counter[5940] = 4'b0000;
    GSharePlugin_logic_mem_counter[5941] = 4'b0000;
    GSharePlugin_logic_mem_counter[5942] = 4'b0000;
    GSharePlugin_logic_mem_counter[5943] = 4'b0000;
    GSharePlugin_logic_mem_counter[5944] = 4'b0000;
    GSharePlugin_logic_mem_counter[5945] = 4'b0000;
    GSharePlugin_logic_mem_counter[5946] = 4'b0000;
    GSharePlugin_logic_mem_counter[5947] = 4'b0000;
    GSharePlugin_logic_mem_counter[5948] = 4'b0000;
    GSharePlugin_logic_mem_counter[5949] = 4'b0000;
    GSharePlugin_logic_mem_counter[5950] = 4'b0000;
    GSharePlugin_logic_mem_counter[5951] = 4'b0000;
    GSharePlugin_logic_mem_counter[5952] = 4'b0000;
    GSharePlugin_logic_mem_counter[5953] = 4'b0000;
    GSharePlugin_logic_mem_counter[5954] = 4'b0000;
    GSharePlugin_logic_mem_counter[5955] = 4'b0000;
    GSharePlugin_logic_mem_counter[5956] = 4'b0000;
    GSharePlugin_logic_mem_counter[5957] = 4'b0000;
    GSharePlugin_logic_mem_counter[5958] = 4'b0000;
    GSharePlugin_logic_mem_counter[5959] = 4'b0000;
    GSharePlugin_logic_mem_counter[5960] = 4'b0000;
    GSharePlugin_logic_mem_counter[5961] = 4'b0000;
    GSharePlugin_logic_mem_counter[5962] = 4'b0000;
    GSharePlugin_logic_mem_counter[5963] = 4'b0000;
    GSharePlugin_logic_mem_counter[5964] = 4'b0000;
    GSharePlugin_logic_mem_counter[5965] = 4'b0000;
    GSharePlugin_logic_mem_counter[5966] = 4'b0000;
    GSharePlugin_logic_mem_counter[5967] = 4'b0000;
    GSharePlugin_logic_mem_counter[5968] = 4'b0000;
    GSharePlugin_logic_mem_counter[5969] = 4'b0000;
    GSharePlugin_logic_mem_counter[5970] = 4'b0000;
    GSharePlugin_logic_mem_counter[5971] = 4'b0000;
    GSharePlugin_logic_mem_counter[5972] = 4'b0000;
    GSharePlugin_logic_mem_counter[5973] = 4'b0000;
    GSharePlugin_logic_mem_counter[5974] = 4'b0000;
    GSharePlugin_logic_mem_counter[5975] = 4'b0000;
    GSharePlugin_logic_mem_counter[5976] = 4'b0000;
    GSharePlugin_logic_mem_counter[5977] = 4'b0000;
    GSharePlugin_logic_mem_counter[5978] = 4'b0000;
    GSharePlugin_logic_mem_counter[5979] = 4'b0000;
    GSharePlugin_logic_mem_counter[5980] = 4'b0000;
    GSharePlugin_logic_mem_counter[5981] = 4'b0000;
    GSharePlugin_logic_mem_counter[5982] = 4'b0000;
    GSharePlugin_logic_mem_counter[5983] = 4'b0000;
    GSharePlugin_logic_mem_counter[5984] = 4'b0000;
    GSharePlugin_logic_mem_counter[5985] = 4'b0000;
    GSharePlugin_logic_mem_counter[5986] = 4'b0000;
    GSharePlugin_logic_mem_counter[5987] = 4'b0000;
    GSharePlugin_logic_mem_counter[5988] = 4'b0000;
    GSharePlugin_logic_mem_counter[5989] = 4'b0000;
    GSharePlugin_logic_mem_counter[5990] = 4'b0000;
    GSharePlugin_logic_mem_counter[5991] = 4'b0000;
    GSharePlugin_logic_mem_counter[5992] = 4'b0000;
    GSharePlugin_logic_mem_counter[5993] = 4'b0000;
    GSharePlugin_logic_mem_counter[5994] = 4'b0000;
    GSharePlugin_logic_mem_counter[5995] = 4'b0000;
    GSharePlugin_logic_mem_counter[5996] = 4'b0000;
    GSharePlugin_logic_mem_counter[5997] = 4'b0000;
    GSharePlugin_logic_mem_counter[5998] = 4'b0000;
    GSharePlugin_logic_mem_counter[5999] = 4'b0000;
    GSharePlugin_logic_mem_counter[6000] = 4'b0000;
    GSharePlugin_logic_mem_counter[6001] = 4'b0000;
    GSharePlugin_logic_mem_counter[6002] = 4'b0000;
    GSharePlugin_logic_mem_counter[6003] = 4'b0000;
    GSharePlugin_logic_mem_counter[6004] = 4'b0000;
    GSharePlugin_logic_mem_counter[6005] = 4'b0000;
    GSharePlugin_logic_mem_counter[6006] = 4'b0000;
    GSharePlugin_logic_mem_counter[6007] = 4'b0000;
    GSharePlugin_logic_mem_counter[6008] = 4'b0000;
    GSharePlugin_logic_mem_counter[6009] = 4'b0000;
    GSharePlugin_logic_mem_counter[6010] = 4'b0000;
    GSharePlugin_logic_mem_counter[6011] = 4'b0000;
    GSharePlugin_logic_mem_counter[6012] = 4'b0000;
    GSharePlugin_logic_mem_counter[6013] = 4'b0000;
    GSharePlugin_logic_mem_counter[6014] = 4'b0000;
    GSharePlugin_logic_mem_counter[6015] = 4'b0000;
    GSharePlugin_logic_mem_counter[6016] = 4'b0000;
    GSharePlugin_logic_mem_counter[6017] = 4'b0000;
    GSharePlugin_logic_mem_counter[6018] = 4'b0000;
    GSharePlugin_logic_mem_counter[6019] = 4'b0000;
    GSharePlugin_logic_mem_counter[6020] = 4'b0000;
    GSharePlugin_logic_mem_counter[6021] = 4'b0000;
    GSharePlugin_logic_mem_counter[6022] = 4'b0000;
    GSharePlugin_logic_mem_counter[6023] = 4'b0000;
    GSharePlugin_logic_mem_counter[6024] = 4'b0000;
    GSharePlugin_logic_mem_counter[6025] = 4'b0000;
    GSharePlugin_logic_mem_counter[6026] = 4'b0000;
    GSharePlugin_logic_mem_counter[6027] = 4'b0000;
    GSharePlugin_logic_mem_counter[6028] = 4'b0000;
    GSharePlugin_logic_mem_counter[6029] = 4'b0000;
    GSharePlugin_logic_mem_counter[6030] = 4'b0000;
    GSharePlugin_logic_mem_counter[6031] = 4'b0000;
    GSharePlugin_logic_mem_counter[6032] = 4'b0000;
    GSharePlugin_logic_mem_counter[6033] = 4'b0000;
    GSharePlugin_logic_mem_counter[6034] = 4'b0000;
    GSharePlugin_logic_mem_counter[6035] = 4'b0000;
    GSharePlugin_logic_mem_counter[6036] = 4'b0000;
    GSharePlugin_logic_mem_counter[6037] = 4'b0000;
    GSharePlugin_logic_mem_counter[6038] = 4'b0000;
    GSharePlugin_logic_mem_counter[6039] = 4'b0000;
    GSharePlugin_logic_mem_counter[6040] = 4'b0000;
    GSharePlugin_logic_mem_counter[6041] = 4'b0000;
    GSharePlugin_logic_mem_counter[6042] = 4'b0000;
    GSharePlugin_logic_mem_counter[6043] = 4'b0000;
    GSharePlugin_logic_mem_counter[6044] = 4'b0000;
    GSharePlugin_logic_mem_counter[6045] = 4'b0000;
    GSharePlugin_logic_mem_counter[6046] = 4'b0000;
    GSharePlugin_logic_mem_counter[6047] = 4'b0000;
    GSharePlugin_logic_mem_counter[6048] = 4'b0000;
    GSharePlugin_logic_mem_counter[6049] = 4'b0000;
    GSharePlugin_logic_mem_counter[6050] = 4'b0000;
    GSharePlugin_logic_mem_counter[6051] = 4'b0000;
    GSharePlugin_logic_mem_counter[6052] = 4'b0000;
    GSharePlugin_logic_mem_counter[6053] = 4'b0000;
    GSharePlugin_logic_mem_counter[6054] = 4'b0000;
    GSharePlugin_logic_mem_counter[6055] = 4'b0000;
    GSharePlugin_logic_mem_counter[6056] = 4'b0000;
    GSharePlugin_logic_mem_counter[6057] = 4'b0000;
    GSharePlugin_logic_mem_counter[6058] = 4'b0000;
    GSharePlugin_logic_mem_counter[6059] = 4'b0000;
    GSharePlugin_logic_mem_counter[6060] = 4'b0000;
    GSharePlugin_logic_mem_counter[6061] = 4'b0000;
    GSharePlugin_logic_mem_counter[6062] = 4'b0000;
    GSharePlugin_logic_mem_counter[6063] = 4'b0000;
    GSharePlugin_logic_mem_counter[6064] = 4'b0000;
    GSharePlugin_logic_mem_counter[6065] = 4'b0000;
    GSharePlugin_logic_mem_counter[6066] = 4'b0000;
    GSharePlugin_logic_mem_counter[6067] = 4'b0000;
    GSharePlugin_logic_mem_counter[6068] = 4'b0000;
    GSharePlugin_logic_mem_counter[6069] = 4'b0000;
    GSharePlugin_logic_mem_counter[6070] = 4'b0000;
    GSharePlugin_logic_mem_counter[6071] = 4'b0000;
    GSharePlugin_logic_mem_counter[6072] = 4'b0000;
    GSharePlugin_logic_mem_counter[6073] = 4'b0000;
    GSharePlugin_logic_mem_counter[6074] = 4'b0000;
    GSharePlugin_logic_mem_counter[6075] = 4'b0000;
    GSharePlugin_logic_mem_counter[6076] = 4'b0000;
    GSharePlugin_logic_mem_counter[6077] = 4'b0000;
    GSharePlugin_logic_mem_counter[6078] = 4'b0000;
    GSharePlugin_logic_mem_counter[6079] = 4'b0000;
    GSharePlugin_logic_mem_counter[6080] = 4'b0000;
    GSharePlugin_logic_mem_counter[6081] = 4'b0000;
    GSharePlugin_logic_mem_counter[6082] = 4'b0000;
    GSharePlugin_logic_mem_counter[6083] = 4'b0000;
    GSharePlugin_logic_mem_counter[6084] = 4'b0000;
    GSharePlugin_logic_mem_counter[6085] = 4'b0000;
    GSharePlugin_logic_mem_counter[6086] = 4'b0000;
    GSharePlugin_logic_mem_counter[6087] = 4'b0000;
    GSharePlugin_logic_mem_counter[6088] = 4'b0000;
    GSharePlugin_logic_mem_counter[6089] = 4'b0000;
    GSharePlugin_logic_mem_counter[6090] = 4'b0000;
    GSharePlugin_logic_mem_counter[6091] = 4'b0000;
    GSharePlugin_logic_mem_counter[6092] = 4'b0000;
    GSharePlugin_logic_mem_counter[6093] = 4'b0000;
    GSharePlugin_logic_mem_counter[6094] = 4'b0000;
    GSharePlugin_logic_mem_counter[6095] = 4'b0000;
    GSharePlugin_logic_mem_counter[6096] = 4'b0000;
    GSharePlugin_logic_mem_counter[6097] = 4'b0000;
    GSharePlugin_logic_mem_counter[6098] = 4'b0000;
    GSharePlugin_logic_mem_counter[6099] = 4'b0000;
    GSharePlugin_logic_mem_counter[6100] = 4'b0000;
    GSharePlugin_logic_mem_counter[6101] = 4'b0000;
    GSharePlugin_logic_mem_counter[6102] = 4'b0000;
    GSharePlugin_logic_mem_counter[6103] = 4'b0000;
    GSharePlugin_logic_mem_counter[6104] = 4'b0000;
    GSharePlugin_logic_mem_counter[6105] = 4'b0000;
    GSharePlugin_logic_mem_counter[6106] = 4'b0000;
    GSharePlugin_logic_mem_counter[6107] = 4'b0000;
    GSharePlugin_logic_mem_counter[6108] = 4'b0000;
    GSharePlugin_logic_mem_counter[6109] = 4'b0000;
    GSharePlugin_logic_mem_counter[6110] = 4'b0000;
    GSharePlugin_logic_mem_counter[6111] = 4'b0000;
    GSharePlugin_logic_mem_counter[6112] = 4'b0000;
    GSharePlugin_logic_mem_counter[6113] = 4'b0000;
    GSharePlugin_logic_mem_counter[6114] = 4'b0000;
    GSharePlugin_logic_mem_counter[6115] = 4'b0000;
    GSharePlugin_logic_mem_counter[6116] = 4'b0000;
    GSharePlugin_logic_mem_counter[6117] = 4'b0000;
    GSharePlugin_logic_mem_counter[6118] = 4'b0000;
    GSharePlugin_logic_mem_counter[6119] = 4'b0000;
    GSharePlugin_logic_mem_counter[6120] = 4'b0000;
    GSharePlugin_logic_mem_counter[6121] = 4'b0000;
    GSharePlugin_logic_mem_counter[6122] = 4'b0000;
    GSharePlugin_logic_mem_counter[6123] = 4'b0000;
    GSharePlugin_logic_mem_counter[6124] = 4'b0000;
    GSharePlugin_logic_mem_counter[6125] = 4'b0000;
    GSharePlugin_logic_mem_counter[6126] = 4'b0000;
    GSharePlugin_logic_mem_counter[6127] = 4'b0000;
    GSharePlugin_logic_mem_counter[6128] = 4'b0000;
    GSharePlugin_logic_mem_counter[6129] = 4'b0000;
    GSharePlugin_logic_mem_counter[6130] = 4'b0000;
    GSharePlugin_logic_mem_counter[6131] = 4'b0000;
    GSharePlugin_logic_mem_counter[6132] = 4'b0000;
    GSharePlugin_logic_mem_counter[6133] = 4'b0000;
    GSharePlugin_logic_mem_counter[6134] = 4'b0000;
    GSharePlugin_logic_mem_counter[6135] = 4'b0000;
    GSharePlugin_logic_mem_counter[6136] = 4'b0000;
    GSharePlugin_logic_mem_counter[6137] = 4'b0000;
    GSharePlugin_logic_mem_counter[6138] = 4'b0000;
    GSharePlugin_logic_mem_counter[6139] = 4'b0000;
    GSharePlugin_logic_mem_counter[6140] = 4'b0000;
    GSharePlugin_logic_mem_counter[6141] = 4'b0000;
    GSharePlugin_logic_mem_counter[6142] = 4'b0000;
    GSharePlugin_logic_mem_counter[6143] = 4'b0000;
    GSharePlugin_logic_mem_counter[6144] = 4'b0000;
    GSharePlugin_logic_mem_counter[6145] = 4'b0000;
    GSharePlugin_logic_mem_counter[6146] = 4'b0000;
    GSharePlugin_logic_mem_counter[6147] = 4'b0000;
    GSharePlugin_logic_mem_counter[6148] = 4'b0000;
    GSharePlugin_logic_mem_counter[6149] = 4'b0000;
    GSharePlugin_logic_mem_counter[6150] = 4'b0000;
    GSharePlugin_logic_mem_counter[6151] = 4'b0000;
    GSharePlugin_logic_mem_counter[6152] = 4'b0000;
    GSharePlugin_logic_mem_counter[6153] = 4'b0000;
    GSharePlugin_logic_mem_counter[6154] = 4'b0000;
    GSharePlugin_logic_mem_counter[6155] = 4'b0000;
    GSharePlugin_logic_mem_counter[6156] = 4'b0000;
    GSharePlugin_logic_mem_counter[6157] = 4'b0000;
    GSharePlugin_logic_mem_counter[6158] = 4'b0000;
    GSharePlugin_logic_mem_counter[6159] = 4'b0000;
    GSharePlugin_logic_mem_counter[6160] = 4'b0000;
    GSharePlugin_logic_mem_counter[6161] = 4'b0000;
    GSharePlugin_logic_mem_counter[6162] = 4'b0000;
    GSharePlugin_logic_mem_counter[6163] = 4'b0000;
    GSharePlugin_logic_mem_counter[6164] = 4'b0000;
    GSharePlugin_logic_mem_counter[6165] = 4'b0000;
    GSharePlugin_logic_mem_counter[6166] = 4'b0000;
    GSharePlugin_logic_mem_counter[6167] = 4'b0000;
    GSharePlugin_logic_mem_counter[6168] = 4'b0000;
    GSharePlugin_logic_mem_counter[6169] = 4'b0000;
    GSharePlugin_logic_mem_counter[6170] = 4'b0000;
    GSharePlugin_logic_mem_counter[6171] = 4'b0000;
    GSharePlugin_logic_mem_counter[6172] = 4'b0000;
    GSharePlugin_logic_mem_counter[6173] = 4'b0000;
    GSharePlugin_logic_mem_counter[6174] = 4'b0000;
    GSharePlugin_logic_mem_counter[6175] = 4'b0000;
    GSharePlugin_logic_mem_counter[6176] = 4'b0000;
    GSharePlugin_logic_mem_counter[6177] = 4'b0000;
    GSharePlugin_logic_mem_counter[6178] = 4'b0000;
    GSharePlugin_logic_mem_counter[6179] = 4'b0000;
    GSharePlugin_logic_mem_counter[6180] = 4'b0000;
    GSharePlugin_logic_mem_counter[6181] = 4'b0000;
    GSharePlugin_logic_mem_counter[6182] = 4'b0000;
    GSharePlugin_logic_mem_counter[6183] = 4'b0000;
    GSharePlugin_logic_mem_counter[6184] = 4'b0000;
    GSharePlugin_logic_mem_counter[6185] = 4'b0000;
    GSharePlugin_logic_mem_counter[6186] = 4'b0000;
    GSharePlugin_logic_mem_counter[6187] = 4'b0000;
    GSharePlugin_logic_mem_counter[6188] = 4'b0000;
    GSharePlugin_logic_mem_counter[6189] = 4'b0000;
    GSharePlugin_logic_mem_counter[6190] = 4'b0000;
    GSharePlugin_logic_mem_counter[6191] = 4'b0000;
    GSharePlugin_logic_mem_counter[6192] = 4'b0000;
    GSharePlugin_logic_mem_counter[6193] = 4'b0000;
    GSharePlugin_logic_mem_counter[6194] = 4'b0000;
    GSharePlugin_logic_mem_counter[6195] = 4'b0000;
    GSharePlugin_logic_mem_counter[6196] = 4'b0000;
    GSharePlugin_logic_mem_counter[6197] = 4'b0000;
    GSharePlugin_logic_mem_counter[6198] = 4'b0000;
    GSharePlugin_logic_mem_counter[6199] = 4'b0000;
    GSharePlugin_logic_mem_counter[6200] = 4'b0000;
    GSharePlugin_logic_mem_counter[6201] = 4'b0000;
    GSharePlugin_logic_mem_counter[6202] = 4'b0000;
    GSharePlugin_logic_mem_counter[6203] = 4'b0000;
    GSharePlugin_logic_mem_counter[6204] = 4'b0000;
    GSharePlugin_logic_mem_counter[6205] = 4'b0000;
    GSharePlugin_logic_mem_counter[6206] = 4'b0000;
    GSharePlugin_logic_mem_counter[6207] = 4'b0000;
    GSharePlugin_logic_mem_counter[6208] = 4'b0000;
    GSharePlugin_logic_mem_counter[6209] = 4'b0000;
    GSharePlugin_logic_mem_counter[6210] = 4'b0000;
    GSharePlugin_logic_mem_counter[6211] = 4'b0000;
    GSharePlugin_logic_mem_counter[6212] = 4'b0000;
    GSharePlugin_logic_mem_counter[6213] = 4'b0000;
    GSharePlugin_logic_mem_counter[6214] = 4'b0000;
    GSharePlugin_logic_mem_counter[6215] = 4'b0000;
    GSharePlugin_logic_mem_counter[6216] = 4'b0000;
    GSharePlugin_logic_mem_counter[6217] = 4'b0000;
    GSharePlugin_logic_mem_counter[6218] = 4'b0000;
    GSharePlugin_logic_mem_counter[6219] = 4'b0000;
    GSharePlugin_logic_mem_counter[6220] = 4'b0000;
    GSharePlugin_logic_mem_counter[6221] = 4'b0000;
    GSharePlugin_logic_mem_counter[6222] = 4'b0000;
    GSharePlugin_logic_mem_counter[6223] = 4'b0000;
    GSharePlugin_logic_mem_counter[6224] = 4'b0000;
    GSharePlugin_logic_mem_counter[6225] = 4'b0000;
    GSharePlugin_logic_mem_counter[6226] = 4'b0000;
    GSharePlugin_logic_mem_counter[6227] = 4'b0000;
    GSharePlugin_logic_mem_counter[6228] = 4'b0000;
    GSharePlugin_logic_mem_counter[6229] = 4'b0000;
    GSharePlugin_logic_mem_counter[6230] = 4'b0000;
    GSharePlugin_logic_mem_counter[6231] = 4'b0000;
    GSharePlugin_logic_mem_counter[6232] = 4'b0000;
    GSharePlugin_logic_mem_counter[6233] = 4'b0000;
    GSharePlugin_logic_mem_counter[6234] = 4'b0000;
    GSharePlugin_logic_mem_counter[6235] = 4'b0000;
    GSharePlugin_logic_mem_counter[6236] = 4'b0000;
    GSharePlugin_logic_mem_counter[6237] = 4'b0000;
    GSharePlugin_logic_mem_counter[6238] = 4'b0000;
    GSharePlugin_logic_mem_counter[6239] = 4'b0000;
    GSharePlugin_logic_mem_counter[6240] = 4'b0000;
    GSharePlugin_logic_mem_counter[6241] = 4'b0000;
    GSharePlugin_logic_mem_counter[6242] = 4'b0000;
    GSharePlugin_logic_mem_counter[6243] = 4'b0000;
    GSharePlugin_logic_mem_counter[6244] = 4'b0000;
    GSharePlugin_logic_mem_counter[6245] = 4'b0000;
    GSharePlugin_logic_mem_counter[6246] = 4'b0000;
    GSharePlugin_logic_mem_counter[6247] = 4'b0000;
    GSharePlugin_logic_mem_counter[6248] = 4'b0000;
    GSharePlugin_logic_mem_counter[6249] = 4'b0000;
    GSharePlugin_logic_mem_counter[6250] = 4'b0000;
    GSharePlugin_logic_mem_counter[6251] = 4'b0000;
    GSharePlugin_logic_mem_counter[6252] = 4'b0000;
    GSharePlugin_logic_mem_counter[6253] = 4'b0000;
    GSharePlugin_logic_mem_counter[6254] = 4'b0000;
    GSharePlugin_logic_mem_counter[6255] = 4'b0000;
    GSharePlugin_logic_mem_counter[6256] = 4'b0000;
    GSharePlugin_logic_mem_counter[6257] = 4'b0000;
    GSharePlugin_logic_mem_counter[6258] = 4'b0000;
    GSharePlugin_logic_mem_counter[6259] = 4'b0000;
    GSharePlugin_logic_mem_counter[6260] = 4'b0000;
    GSharePlugin_logic_mem_counter[6261] = 4'b0000;
    GSharePlugin_logic_mem_counter[6262] = 4'b0000;
    GSharePlugin_logic_mem_counter[6263] = 4'b0000;
    GSharePlugin_logic_mem_counter[6264] = 4'b0000;
    GSharePlugin_logic_mem_counter[6265] = 4'b0000;
    GSharePlugin_logic_mem_counter[6266] = 4'b0000;
    GSharePlugin_logic_mem_counter[6267] = 4'b0000;
    GSharePlugin_logic_mem_counter[6268] = 4'b0000;
    GSharePlugin_logic_mem_counter[6269] = 4'b0000;
    GSharePlugin_logic_mem_counter[6270] = 4'b0000;
    GSharePlugin_logic_mem_counter[6271] = 4'b0000;
    GSharePlugin_logic_mem_counter[6272] = 4'b0000;
    GSharePlugin_logic_mem_counter[6273] = 4'b0000;
    GSharePlugin_logic_mem_counter[6274] = 4'b0000;
    GSharePlugin_logic_mem_counter[6275] = 4'b0000;
    GSharePlugin_logic_mem_counter[6276] = 4'b0000;
    GSharePlugin_logic_mem_counter[6277] = 4'b0000;
    GSharePlugin_logic_mem_counter[6278] = 4'b0000;
    GSharePlugin_logic_mem_counter[6279] = 4'b0000;
    GSharePlugin_logic_mem_counter[6280] = 4'b0000;
    GSharePlugin_logic_mem_counter[6281] = 4'b0000;
    GSharePlugin_logic_mem_counter[6282] = 4'b0000;
    GSharePlugin_logic_mem_counter[6283] = 4'b0000;
    GSharePlugin_logic_mem_counter[6284] = 4'b0000;
    GSharePlugin_logic_mem_counter[6285] = 4'b0000;
    GSharePlugin_logic_mem_counter[6286] = 4'b0000;
    GSharePlugin_logic_mem_counter[6287] = 4'b0000;
    GSharePlugin_logic_mem_counter[6288] = 4'b0000;
    GSharePlugin_logic_mem_counter[6289] = 4'b0000;
    GSharePlugin_logic_mem_counter[6290] = 4'b0000;
    GSharePlugin_logic_mem_counter[6291] = 4'b0000;
    GSharePlugin_logic_mem_counter[6292] = 4'b0000;
    GSharePlugin_logic_mem_counter[6293] = 4'b0000;
    GSharePlugin_logic_mem_counter[6294] = 4'b0000;
    GSharePlugin_logic_mem_counter[6295] = 4'b0000;
    GSharePlugin_logic_mem_counter[6296] = 4'b0000;
    GSharePlugin_logic_mem_counter[6297] = 4'b0000;
    GSharePlugin_logic_mem_counter[6298] = 4'b0000;
    GSharePlugin_logic_mem_counter[6299] = 4'b0000;
    GSharePlugin_logic_mem_counter[6300] = 4'b0000;
    GSharePlugin_logic_mem_counter[6301] = 4'b0000;
    GSharePlugin_logic_mem_counter[6302] = 4'b0000;
    GSharePlugin_logic_mem_counter[6303] = 4'b0000;
    GSharePlugin_logic_mem_counter[6304] = 4'b0000;
    GSharePlugin_logic_mem_counter[6305] = 4'b0000;
    GSharePlugin_logic_mem_counter[6306] = 4'b0000;
    GSharePlugin_logic_mem_counter[6307] = 4'b0000;
    GSharePlugin_logic_mem_counter[6308] = 4'b0000;
    GSharePlugin_logic_mem_counter[6309] = 4'b0000;
    GSharePlugin_logic_mem_counter[6310] = 4'b0000;
    GSharePlugin_logic_mem_counter[6311] = 4'b0000;
    GSharePlugin_logic_mem_counter[6312] = 4'b0000;
    GSharePlugin_logic_mem_counter[6313] = 4'b0000;
    GSharePlugin_logic_mem_counter[6314] = 4'b0000;
    GSharePlugin_logic_mem_counter[6315] = 4'b0000;
    GSharePlugin_logic_mem_counter[6316] = 4'b0000;
    GSharePlugin_logic_mem_counter[6317] = 4'b0000;
    GSharePlugin_logic_mem_counter[6318] = 4'b0000;
    GSharePlugin_logic_mem_counter[6319] = 4'b0000;
    GSharePlugin_logic_mem_counter[6320] = 4'b0000;
    GSharePlugin_logic_mem_counter[6321] = 4'b0000;
    GSharePlugin_logic_mem_counter[6322] = 4'b0000;
    GSharePlugin_logic_mem_counter[6323] = 4'b0000;
    GSharePlugin_logic_mem_counter[6324] = 4'b0000;
    GSharePlugin_logic_mem_counter[6325] = 4'b0000;
    GSharePlugin_logic_mem_counter[6326] = 4'b0000;
    GSharePlugin_logic_mem_counter[6327] = 4'b0000;
    GSharePlugin_logic_mem_counter[6328] = 4'b0000;
    GSharePlugin_logic_mem_counter[6329] = 4'b0000;
    GSharePlugin_logic_mem_counter[6330] = 4'b0000;
    GSharePlugin_logic_mem_counter[6331] = 4'b0000;
    GSharePlugin_logic_mem_counter[6332] = 4'b0000;
    GSharePlugin_logic_mem_counter[6333] = 4'b0000;
    GSharePlugin_logic_mem_counter[6334] = 4'b0000;
    GSharePlugin_logic_mem_counter[6335] = 4'b0000;
    GSharePlugin_logic_mem_counter[6336] = 4'b0000;
    GSharePlugin_logic_mem_counter[6337] = 4'b0000;
    GSharePlugin_logic_mem_counter[6338] = 4'b0000;
    GSharePlugin_logic_mem_counter[6339] = 4'b0000;
    GSharePlugin_logic_mem_counter[6340] = 4'b0000;
    GSharePlugin_logic_mem_counter[6341] = 4'b0000;
    GSharePlugin_logic_mem_counter[6342] = 4'b0000;
    GSharePlugin_logic_mem_counter[6343] = 4'b0000;
    GSharePlugin_logic_mem_counter[6344] = 4'b0000;
    GSharePlugin_logic_mem_counter[6345] = 4'b0000;
    GSharePlugin_logic_mem_counter[6346] = 4'b0000;
    GSharePlugin_logic_mem_counter[6347] = 4'b0000;
    GSharePlugin_logic_mem_counter[6348] = 4'b0000;
    GSharePlugin_logic_mem_counter[6349] = 4'b0000;
    GSharePlugin_logic_mem_counter[6350] = 4'b0000;
    GSharePlugin_logic_mem_counter[6351] = 4'b0000;
    GSharePlugin_logic_mem_counter[6352] = 4'b0000;
    GSharePlugin_logic_mem_counter[6353] = 4'b0000;
    GSharePlugin_logic_mem_counter[6354] = 4'b0000;
    GSharePlugin_logic_mem_counter[6355] = 4'b0000;
    GSharePlugin_logic_mem_counter[6356] = 4'b0000;
    GSharePlugin_logic_mem_counter[6357] = 4'b0000;
    GSharePlugin_logic_mem_counter[6358] = 4'b0000;
    GSharePlugin_logic_mem_counter[6359] = 4'b0000;
    GSharePlugin_logic_mem_counter[6360] = 4'b0000;
    GSharePlugin_logic_mem_counter[6361] = 4'b0000;
    GSharePlugin_logic_mem_counter[6362] = 4'b0000;
    GSharePlugin_logic_mem_counter[6363] = 4'b0000;
    GSharePlugin_logic_mem_counter[6364] = 4'b0000;
    GSharePlugin_logic_mem_counter[6365] = 4'b0000;
    GSharePlugin_logic_mem_counter[6366] = 4'b0000;
    GSharePlugin_logic_mem_counter[6367] = 4'b0000;
    GSharePlugin_logic_mem_counter[6368] = 4'b0000;
    GSharePlugin_logic_mem_counter[6369] = 4'b0000;
    GSharePlugin_logic_mem_counter[6370] = 4'b0000;
    GSharePlugin_logic_mem_counter[6371] = 4'b0000;
    GSharePlugin_logic_mem_counter[6372] = 4'b0000;
    GSharePlugin_logic_mem_counter[6373] = 4'b0000;
    GSharePlugin_logic_mem_counter[6374] = 4'b0000;
    GSharePlugin_logic_mem_counter[6375] = 4'b0000;
    GSharePlugin_logic_mem_counter[6376] = 4'b0000;
    GSharePlugin_logic_mem_counter[6377] = 4'b0000;
    GSharePlugin_logic_mem_counter[6378] = 4'b0000;
    GSharePlugin_logic_mem_counter[6379] = 4'b0000;
    GSharePlugin_logic_mem_counter[6380] = 4'b0000;
    GSharePlugin_logic_mem_counter[6381] = 4'b0000;
    GSharePlugin_logic_mem_counter[6382] = 4'b0000;
    GSharePlugin_logic_mem_counter[6383] = 4'b0000;
    GSharePlugin_logic_mem_counter[6384] = 4'b0000;
    GSharePlugin_logic_mem_counter[6385] = 4'b0000;
    GSharePlugin_logic_mem_counter[6386] = 4'b0000;
    GSharePlugin_logic_mem_counter[6387] = 4'b0000;
    GSharePlugin_logic_mem_counter[6388] = 4'b0000;
    GSharePlugin_logic_mem_counter[6389] = 4'b0000;
    GSharePlugin_logic_mem_counter[6390] = 4'b0000;
    GSharePlugin_logic_mem_counter[6391] = 4'b0000;
    GSharePlugin_logic_mem_counter[6392] = 4'b0000;
    GSharePlugin_logic_mem_counter[6393] = 4'b0000;
    GSharePlugin_logic_mem_counter[6394] = 4'b0000;
    GSharePlugin_logic_mem_counter[6395] = 4'b0000;
    GSharePlugin_logic_mem_counter[6396] = 4'b0000;
    GSharePlugin_logic_mem_counter[6397] = 4'b0000;
    GSharePlugin_logic_mem_counter[6398] = 4'b0000;
    GSharePlugin_logic_mem_counter[6399] = 4'b0000;
    GSharePlugin_logic_mem_counter[6400] = 4'b0000;
    GSharePlugin_logic_mem_counter[6401] = 4'b0000;
    GSharePlugin_logic_mem_counter[6402] = 4'b0000;
    GSharePlugin_logic_mem_counter[6403] = 4'b0000;
    GSharePlugin_logic_mem_counter[6404] = 4'b0000;
    GSharePlugin_logic_mem_counter[6405] = 4'b0000;
    GSharePlugin_logic_mem_counter[6406] = 4'b0000;
    GSharePlugin_logic_mem_counter[6407] = 4'b0000;
    GSharePlugin_logic_mem_counter[6408] = 4'b0000;
    GSharePlugin_logic_mem_counter[6409] = 4'b0000;
    GSharePlugin_logic_mem_counter[6410] = 4'b0000;
    GSharePlugin_logic_mem_counter[6411] = 4'b0000;
    GSharePlugin_logic_mem_counter[6412] = 4'b0000;
    GSharePlugin_logic_mem_counter[6413] = 4'b0000;
    GSharePlugin_logic_mem_counter[6414] = 4'b0000;
    GSharePlugin_logic_mem_counter[6415] = 4'b0000;
    GSharePlugin_logic_mem_counter[6416] = 4'b0000;
    GSharePlugin_logic_mem_counter[6417] = 4'b0000;
    GSharePlugin_logic_mem_counter[6418] = 4'b0000;
    GSharePlugin_logic_mem_counter[6419] = 4'b0000;
    GSharePlugin_logic_mem_counter[6420] = 4'b0000;
    GSharePlugin_logic_mem_counter[6421] = 4'b0000;
    GSharePlugin_logic_mem_counter[6422] = 4'b0000;
    GSharePlugin_logic_mem_counter[6423] = 4'b0000;
    GSharePlugin_logic_mem_counter[6424] = 4'b0000;
    GSharePlugin_logic_mem_counter[6425] = 4'b0000;
    GSharePlugin_logic_mem_counter[6426] = 4'b0000;
    GSharePlugin_logic_mem_counter[6427] = 4'b0000;
    GSharePlugin_logic_mem_counter[6428] = 4'b0000;
    GSharePlugin_logic_mem_counter[6429] = 4'b0000;
    GSharePlugin_logic_mem_counter[6430] = 4'b0000;
    GSharePlugin_logic_mem_counter[6431] = 4'b0000;
    GSharePlugin_logic_mem_counter[6432] = 4'b0000;
    GSharePlugin_logic_mem_counter[6433] = 4'b0000;
    GSharePlugin_logic_mem_counter[6434] = 4'b0000;
    GSharePlugin_logic_mem_counter[6435] = 4'b0000;
    GSharePlugin_logic_mem_counter[6436] = 4'b0000;
    GSharePlugin_logic_mem_counter[6437] = 4'b0000;
    GSharePlugin_logic_mem_counter[6438] = 4'b0000;
    GSharePlugin_logic_mem_counter[6439] = 4'b0000;
    GSharePlugin_logic_mem_counter[6440] = 4'b0000;
    GSharePlugin_logic_mem_counter[6441] = 4'b0000;
    GSharePlugin_logic_mem_counter[6442] = 4'b0000;
    GSharePlugin_logic_mem_counter[6443] = 4'b0000;
    GSharePlugin_logic_mem_counter[6444] = 4'b0000;
    GSharePlugin_logic_mem_counter[6445] = 4'b0000;
    GSharePlugin_logic_mem_counter[6446] = 4'b0000;
    GSharePlugin_logic_mem_counter[6447] = 4'b0000;
    GSharePlugin_logic_mem_counter[6448] = 4'b0000;
    GSharePlugin_logic_mem_counter[6449] = 4'b0000;
    GSharePlugin_logic_mem_counter[6450] = 4'b0000;
    GSharePlugin_logic_mem_counter[6451] = 4'b0000;
    GSharePlugin_logic_mem_counter[6452] = 4'b0000;
    GSharePlugin_logic_mem_counter[6453] = 4'b0000;
    GSharePlugin_logic_mem_counter[6454] = 4'b0000;
    GSharePlugin_logic_mem_counter[6455] = 4'b0000;
    GSharePlugin_logic_mem_counter[6456] = 4'b0000;
    GSharePlugin_logic_mem_counter[6457] = 4'b0000;
    GSharePlugin_logic_mem_counter[6458] = 4'b0000;
    GSharePlugin_logic_mem_counter[6459] = 4'b0000;
    GSharePlugin_logic_mem_counter[6460] = 4'b0000;
    GSharePlugin_logic_mem_counter[6461] = 4'b0000;
    GSharePlugin_logic_mem_counter[6462] = 4'b0000;
    GSharePlugin_logic_mem_counter[6463] = 4'b0000;
    GSharePlugin_logic_mem_counter[6464] = 4'b0000;
    GSharePlugin_logic_mem_counter[6465] = 4'b0000;
    GSharePlugin_logic_mem_counter[6466] = 4'b0000;
    GSharePlugin_logic_mem_counter[6467] = 4'b0000;
    GSharePlugin_logic_mem_counter[6468] = 4'b0000;
    GSharePlugin_logic_mem_counter[6469] = 4'b0000;
    GSharePlugin_logic_mem_counter[6470] = 4'b0000;
    GSharePlugin_logic_mem_counter[6471] = 4'b0000;
    GSharePlugin_logic_mem_counter[6472] = 4'b0000;
    GSharePlugin_logic_mem_counter[6473] = 4'b0000;
    GSharePlugin_logic_mem_counter[6474] = 4'b0000;
    GSharePlugin_logic_mem_counter[6475] = 4'b0000;
    GSharePlugin_logic_mem_counter[6476] = 4'b0000;
    GSharePlugin_logic_mem_counter[6477] = 4'b0000;
    GSharePlugin_logic_mem_counter[6478] = 4'b0000;
    GSharePlugin_logic_mem_counter[6479] = 4'b0000;
    GSharePlugin_logic_mem_counter[6480] = 4'b0000;
    GSharePlugin_logic_mem_counter[6481] = 4'b0000;
    GSharePlugin_logic_mem_counter[6482] = 4'b0000;
    GSharePlugin_logic_mem_counter[6483] = 4'b0000;
    GSharePlugin_logic_mem_counter[6484] = 4'b0000;
    GSharePlugin_logic_mem_counter[6485] = 4'b0000;
    GSharePlugin_logic_mem_counter[6486] = 4'b0000;
    GSharePlugin_logic_mem_counter[6487] = 4'b0000;
    GSharePlugin_logic_mem_counter[6488] = 4'b0000;
    GSharePlugin_logic_mem_counter[6489] = 4'b0000;
    GSharePlugin_logic_mem_counter[6490] = 4'b0000;
    GSharePlugin_logic_mem_counter[6491] = 4'b0000;
    GSharePlugin_logic_mem_counter[6492] = 4'b0000;
    GSharePlugin_logic_mem_counter[6493] = 4'b0000;
    GSharePlugin_logic_mem_counter[6494] = 4'b0000;
    GSharePlugin_logic_mem_counter[6495] = 4'b0000;
    GSharePlugin_logic_mem_counter[6496] = 4'b0000;
    GSharePlugin_logic_mem_counter[6497] = 4'b0000;
    GSharePlugin_logic_mem_counter[6498] = 4'b0000;
    GSharePlugin_logic_mem_counter[6499] = 4'b0000;
    GSharePlugin_logic_mem_counter[6500] = 4'b0000;
    GSharePlugin_logic_mem_counter[6501] = 4'b0000;
    GSharePlugin_logic_mem_counter[6502] = 4'b0000;
    GSharePlugin_logic_mem_counter[6503] = 4'b0000;
    GSharePlugin_logic_mem_counter[6504] = 4'b0000;
    GSharePlugin_logic_mem_counter[6505] = 4'b0000;
    GSharePlugin_logic_mem_counter[6506] = 4'b0000;
    GSharePlugin_logic_mem_counter[6507] = 4'b0000;
    GSharePlugin_logic_mem_counter[6508] = 4'b0000;
    GSharePlugin_logic_mem_counter[6509] = 4'b0000;
    GSharePlugin_logic_mem_counter[6510] = 4'b0000;
    GSharePlugin_logic_mem_counter[6511] = 4'b0000;
    GSharePlugin_logic_mem_counter[6512] = 4'b0000;
    GSharePlugin_logic_mem_counter[6513] = 4'b0000;
    GSharePlugin_logic_mem_counter[6514] = 4'b0000;
    GSharePlugin_logic_mem_counter[6515] = 4'b0000;
    GSharePlugin_logic_mem_counter[6516] = 4'b0000;
    GSharePlugin_logic_mem_counter[6517] = 4'b0000;
    GSharePlugin_logic_mem_counter[6518] = 4'b0000;
    GSharePlugin_logic_mem_counter[6519] = 4'b0000;
    GSharePlugin_logic_mem_counter[6520] = 4'b0000;
    GSharePlugin_logic_mem_counter[6521] = 4'b0000;
    GSharePlugin_logic_mem_counter[6522] = 4'b0000;
    GSharePlugin_logic_mem_counter[6523] = 4'b0000;
    GSharePlugin_logic_mem_counter[6524] = 4'b0000;
    GSharePlugin_logic_mem_counter[6525] = 4'b0000;
    GSharePlugin_logic_mem_counter[6526] = 4'b0000;
    GSharePlugin_logic_mem_counter[6527] = 4'b0000;
    GSharePlugin_logic_mem_counter[6528] = 4'b0000;
    GSharePlugin_logic_mem_counter[6529] = 4'b0000;
    GSharePlugin_logic_mem_counter[6530] = 4'b0000;
    GSharePlugin_logic_mem_counter[6531] = 4'b0000;
    GSharePlugin_logic_mem_counter[6532] = 4'b0000;
    GSharePlugin_logic_mem_counter[6533] = 4'b0000;
    GSharePlugin_logic_mem_counter[6534] = 4'b0000;
    GSharePlugin_logic_mem_counter[6535] = 4'b0000;
    GSharePlugin_logic_mem_counter[6536] = 4'b0000;
    GSharePlugin_logic_mem_counter[6537] = 4'b0000;
    GSharePlugin_logic_mem_counter[6538] = 4'b0000;
    GSharePlugin_logic_mem_counter[6539] = 4'b0000;
    GSharePlugin_logic_mem_counter[6540] = 4'b0000;
    GSharePlugin_logic_mem_counter[6541] = 4'b0000;
    GSharePlugin_logic_mem_counter[6542] = 4'b0000;
    GSharePlugin_logic_mem_counter[6543] = 4'b0000;
    GSharePlugin_logic_mem_counter[6544] = 4'b0000;
    GSharePlugin_logic_mem_counter[6545] = 4'b0000;
    GSharePlugin_logic_mem_counter[6546] = 4'b0000;
    GSharePlugin_logic_mem_counter[6547] = 4'b0000;
    GSharePlugin_logic_mem_counter[6548] = 4'b0000;
    GSharePlugin_logic_mem_counter[6549] = 4'b0000;
    GSharePlugin_logic_mem_counter[6550] = 4'b0000;
    GSharePlugin_logic_mem_counter[6551] = 4'b0000;
    GSharePlugin_logic_mem_counter[6552] = 4'b0000;
    GSharePlugin_logic_mem_counter[6553] = 4'b0000;
    GSharePlugin_logic_mem_counter[6554] = 4'b0000;
    GSharePlugin_logic_mem_counter[6555] = 4'b0000;
    GSharePlugin_logic_mem_counter[6556] = 4'b0000;
    GSharePlugin_logic_mem_counter[6557] = 4'b0000;
    GSharePlugin_logic_mem_counter[6558] = 4'b0000;
    GSharePlugin_logic_mem_counter[6559] = 4'b0000;
    GSharePlugin_logic_mem_counter[6560] = 4'b0000;
    GSharePlugin_logic_mem_counter[6561] = 4'b0000;
    GSharePlugin_logic_mem_counter[6562] = 4'b0000;
    GSharePlugin_logic_mem_counter[6563] = 4'b0000;
    GSharePlugin_logic_mem_counter[6564] = 4'b0000;
    GSharePlugin_logic_mem_counter[6565] = 4'b0000;
    GSharePlugin_logic_mem_counter[6566] = 4'b0000;
    GSharePlugin_logic_mem_counter[6567] = 4'b0000;
    GSharePlugin_logic_mem_counter[6568] = 4'b0000;
    GSharePlugin_logic_mem_counter[6569] = 4'b0000;
    GSharePlugin_logic_mem_counter[6570] = 4'b0000;
    GSharePlugin_logic_mem_counter[6571] = 4'b0000;
    GSharePlugin_logic_mem_counter[6572] = 4'b0000;
    GSharePlugin_logic_mem_counter[6573] = 4'b0000;
    GSharePlugin_logic_mem_counter[6574] = 4'b0000;
    GSharePlugin_logic_mem_counter[6575] = 4'b0000;
    GSharePlugin_logic_mem_counter[6576] = 4'b0000;
    GSharePlugin_logic_mem_counter[6577] = 4'b0000;
    GSharePlugin_logic_mem_counter[6578] = 4'b0000;
    GSharePlugin_logic_mem_counter[6579] = 4'b0000;
    GSharePlugin_logic_mem_counter[6580] = 4'b0000;
    GSharePlugin_logic_mem_counter[6581] = 4'b0000;
    GSharePlugin_logic_mem_counter[6582] = 4'b0000;
    GSharePlugin_logic_mem_counter[6583] = 4'b0000;
    GSharePlugin_logic_mem_counter[6584] = 4'b0000;
    GSharePlugin_logic_mem_counter[6585] = 4'b0000;
    GSharePlugin_logic_mem_counter[6586] = 4'b0000;
    GSharePlugin_logic_mem_counter[6587] = 4'b0000;
    GSharePlugin_logic_mem_counter[6588] = 4'b0000;
    GSharePlugin_logic_mem_counter[6589] = 4'b0000;
    GSharePlugin_logic_mem_counter[6590] = 4'b0000;
    GSharePlugin_logic_mem_counter[6591] = 4'b0000;
    GSharePlugin_logic_mem_counter[6592] = 4'b0000;
    GSharePlugin_logic_mem_counter[6593] = 4'b0000;
    GSharePlugin_logic_mem_counter[6594] = 4'b0000;
    GSharePlugin_logic_mem_counter[6595] = 4'b0000;
    GSharePlugin_logic_mem_counter[6596] = 4'b0000;
    GSharePlugin_logic_mem_counter[6597] = 4'b0000;
    GSharePlugin_logic_mem_counter[6598] = 4'b0000;
    GSharePlugin_logic_mem_counter[6599] = 4'b0000;
    GSharePlugin_logic_mem_counter[6600] = 4'b0000;
    GSharePlugin_logic_mem_counter[6601] = 4'b0000;
    GSharePlugin_logic_mem_counter[6602] = 4'b0000;
    GSharePlugin_logic_mem_counter[6603] = 4'b0000;
    GSharePlugin_logic_mem_counter[6604] = 4'b0000;
    GSharePlugin_logic_mem_counter[6605] = 4'b0000;
    GSharePlugin_logic_mem_counter[6606] = 4'b0000;
    GSharePlugin_logic_mem_counter[6607] = 4'b0000;
    GSharePlugin_logic_mem_counter[6608] = 4'b0000;
    GSharePlugin_logic_mem_counter[6609] = 4'b0000;
    GSharePlugin_logic_mem_counter[6610] = 4'b0000;
    GSharePlugin_logic_mem_counter[6611] = 4'b0000;
    GSharePlugin_logic_mem_counter[6612] = 4'b0000;
    GSharePlugin_logic_mem_counter[6613] = 4'b0000;
    GSharePlugin_logic_mem_counter[6614] = 4'b0000;
    GSharePlugin_logic_mem_counter[6615] = 4'b0000;
    GSharePlugin_logic_mem_counter[6616] = 4'b0000;
    GSharePlugin_logic_mem_counter[6617] = 4'b0000;
    GSharePlugin_logic_mem_counter[6618] = 4'b0000;
    GSharePlugin_logic_mem_counter[6619] = 4'b0000;
    GSharePlugin_logic_mem_counter[6620] = 4'b0000;
    GSharePlugin_logic_mem_counter[6621] = 4'b0000;
    GSharePlugin_logic_mem_counter[6622] = 4'b0000;
    GSharePlugin_logic_mem_counter[6623] = 4'b0000;
    GSharePlugin_logic_mem_counter[6624] = 4'b0000;
    GSharePlugin_logic_mem_counter[6625] = 4'b0000;
    GSharePlugin_logic_mem_counter[6626] = 4'b0000;
    GSharePlugin_logic_mem_counter[6627] = 4'b0000;
    GSharePlugin_logic_mem_counter[6628] = 4'b0000;
    GSharePlugin_logic_mem_counter[6629] = 4'b0000;
    GSharePlugin_logic_mem_counter[6630] = 4'b0000;
    GSharePlugin_logic_mem_counter[6631] = 4'b0000;
    GSharePlugin_logic_mem_counter[6632] = 4'b0000;
    GSharePlugin_logic_mem_counter[6633] = 4'b0000;
    GSharePlugin_logic_mem_counter[6634] = 4'b0000;
    GSharePlugin_logic_mem_counter[6635] = 4'b0000;
    GSharePlugin_logic_mem_counter[6636] = 4'b0000;
    GSharePlugin_logic_mem_counter[6637] = 4'b0000;
    GSharePlugin_logic_mem_counter[6638] = 4'b0000;
    GSharePlugin_logic_mem_counter[6639] = 4'b0000;
    GSharePlugin_logic_mem_counter[6640] = 4'b0000;
    GSharePlugin_logic_mem_counter[6641] = 4'b0000;
    GSharePlugin_logic_mem_counter[6642] = 4'b0000;
    GSharePlugin_logic_mem_counter[6643] = 4'b0000;
    GSharePlugin_logic_mem_counter[6644] = 4'b0000;
    GSharePlugin_logic_mem_counter[6645] = 4'b0000;
    GSharePlugin_logic_mem_counter[6646] = 4'b0000;
    GSharePlugin_logic_mem_counter[6647] = 4'b0000;
    GSharePlugin_logic_mem_counter[6648] = 4'b0000;
    GSharePlugin_logic_mem_counter[6649] = 4'b0000;
    GSharePlugin_logic_mem_counter[6650] = 4'b0000;
    GSharePlugin_logic_mem_counter[6651] = 4'b0000;
    GSharePlugin_logic_mem_counter[6652] = 4'b0000;
    GSharePlugin_logic_mem_counter[6653] = 4'b0000;
    GSharePlugin_logic_mem_counter[6654] = 4'b0000;
    GSharePlugin_logic_mem_counter[6655] = 4'b0000;
    GSharePlugin_logic_mem_counter[6656] = 4'b0000;
    GSharePlugin_logic_mem_counter[6657] = 4'b0000;
    GSharePlugin_logic_mem_counter[6658] = 4'b0000;
    GSharePlugin_logic_mem_counter[6659] = 4'b0000;
    GSharePlugin_logic_mem_counter[6660] = 4'b0000;
    GSharePlugin_logic_mem_counter[6661] = 4'b0000;
    GSharePlugin_logic_mem_counter[6662] = 4'b0000;
    GSharePlugin_logic_mem_counter[6663] = 4'b0000;
    GSharePlugin_logic_mem_counter[6664] = 4'b0000;
    GSharePlugin_logic_mem_counter[6665] = 4'b0000;
    GSharePlugin_logic_mem_counter[6666] = 4'b0000;
    GSharePlugin_logic_mem_counter[6667] = 4'b0000;
    GSharePlugin_logic_mem_counter[6668] = 4'b0000;
    GSharePlugin_logic_mem_counter[6669] = 4'b0000;
    GSharePlugin_logic_mem_counter[6670] = 4'b0000;
    GSharePlugin_logic_mem_counter[6671] = 4'b0000;
    GSharePlugin_logic_mem_counter[6672] = 4'b0000;
    GSharePlugin_logic_mem_counter[6673] = 4'b0000;
    GSharePlugin_logic_mem_counter[6674] = 4'b0000;
    GSharePlugin_logic_mem_counter[6675] = 4'b0000;
    GSharePlugin_logic_mem_counter[6676] = 4'b0000;
    GSharePlugin_logic_mem_counter[6677] = 4'b0000;
    GSharePlugin_logic_mem_counter[6678] = 4'b0000;
    GSharePlugin_logic_mem_counter[6679] = 4'b0000;
    GSharePlugin_logic_mem_counter[6680] = 4'b0000;
    GSharePlugin_logic_mem_counter[6681] = 4'b0000;
    GSharePlugin_logic_mem_counter[6682] = 4'b0000;
    GSharePlugin_logic_mem_counter[6683] = 4'b0000;
    GSharePlugin_logic_mem_counter[6684] = 4'b0000;
    GSharePlugin_logic_mem_counter[6685] = 4'b0000;
    GSharePlugin_logic_mem_counter[6686] = 4'b0000;
    GSharePlugin_logic_mem_counter[6687] = 4'b0000;
    GSharePlugin_logic_mem_counter[6688] = 4'b0000;
    GSharePlugin_logic_mem_counter[6689] = 4'b0000;
    GSharePlugin_logic_mem_counter[6690] = 4'b0000;
    GSharePlugin_logic_mem_counter[6691] = 4'b0000;
    GSharePlugin_logic_mem_counter[6692] = 4'b0000;
    GSharePlugin_logic_mem_counter[6693] = 4'b0000;
    GSharePlugin_logic_mem_counter[6694] = 4'b0000;
    GSharePlugin_logic_mem_counter[6695] = 4'b0000;
    GSharePlugin_logic_mem_counter[6696] = 4'b0000;
    GSharePlugin_logic_mem_counter[6697] = 4'b0000;
    GSharePlugin_logic_mem_counter[6698] = 4'b0000;
    GSharePlugin_logic_mem_counter[6699] = 4'b0000;
    GSharePlugin_logic_mem_counter[6700] = 4'b0000;
    GSharePlugin_logic_mem_counter[6701] = 4'b0000;
    GSharePlugin_logic_mem_counter[6702] = 4'b0000;
    GSharePlugin_logic_mem_counter[6703] = 4'b0000;
    GSharePlugin_logic_mem_counter[6704] = 4'b0000;
    GSharePlugin_logic_mem_counter[6705] = 4'b0000;
    GSharePlugin_logic_mem_counter[6706] = 4'b0000;
    GSharePlugin_logic_mem_counter[6707] = 4'b0000;
    GSharePlugin_logic_mem_counter[6708] = 4'b0000;
    GSharePlugin_logic_mem_counter[6709] = 4'b0000;
    GSharePlugin_logic_mem_counter[6710] = 4'b0000;
    GSharePlugin_logic_mem_counter[6711] = 4'b0000;
    GSharePlugin_logic_mem_counter[6712] = 4'b0000;
    GSharePlugin_logic_mem_counter[6713] = 4'b0000;
    GSharePlugin_logic_mem_counter[6714] = 4'b0000;
    GSharePlugin_logic_mem_counter[6715] = 4'b0000;
    GSharePlugin_logic_mem_counter[6716] = 4'b0000;
    GSharePlugin_logic_mem_counter[6717] = 4'b0000;
    GSharePlugin_logic_mem_counter[6718] = 4'b0000;
    GSharePlugin_logic_mem_counter[6719] = 4'b0000;
    GSharePlugin_logic_mem_counter[6720] = 4'b0000;
    GSharePlugin_logic_mem_counter[6721] = 4'b0000;
    GSharePlugin_logic_mem_counter[6722] = 4'b0000;
    GSharePlugin_logic_mem_counter[6723] = 4'b0000;
    GSharePlugin_logic_mem_counter[6724] = 4'b0000;
    GSharePlugin_logic_mem_counter[6725] = 4'b0000;
    GSharePlugin_logic_mem_counter[6726] = 4'b0000;
    GSharePlugin_logic_mem_counter[6727] = 4'b0000;
    GSharePlugin_logic_mem_counter[6728] = 4'b0000;
    GSharePlugin_logic_mem_counter[6729] = 4'b0000;
    GSharePlugin_logic_mem_counter[6730] = 4'b0000;
    GSharePlugin_logic_mem_counter[6731] = 4'b0000;
    GSharePlugin_logic_mem_counter[6732] = 4'b0000;
    GSharePlugin_logic_mem_counter[6733] = 4'b0000;
    GSharePlugin_logic_mem_counter[6734] = 4'b0000;
    GSharePlugin_logic_mem_counter[6735] = 4'b0000;
    GSharePlugin_logic_mem_counter[6736] = 4'b0000;
    GSharePlugin_logic_mem_counter[6737] = 4'b0000;
    GSharePlugin_logic_mem_counter[6738] = 4'b0000;
    GSharePlugin_logic_mem_counter[6739] = 4'b0000;
    GSharePlugin_logic_mem_counter[6740] = 4'b0000;
    GSharePlugin_logic_mem_counter[6741] = 4'b0000;
    GSharePlugin_logic_mem_counter[6742] = 4'b0000;
    GSharePlugin_logic_mem_counter[6743] = 4'b0000;
    GSharePlugin_logic_mem_counter[6744] = 4'b0000;
    GSharePlugin_logic_mem_counter[6745] = 4'b0000;
    GSharePlugin_logic_mem_counter[6746] = 4'b0000;
    GSharePlugin_logic_mem_counter[6747] = 4'b0000;
    GSharePlugin_logic_mem_counter[6748] = 4'b0000;
    GSharePlugin_logic_mem_counter[6749] = 4'b0000;
    GSharePlugin_logic_mem_counter[6750] = 4'b0000;
    GSharePlugin_logic_mem_counter[6751] = 4'b0000;
    GSharePlugin_logic_mem_counter[6752] = 4'b0000;
    GSharePlugin_logic_mem_counter[6753] = 4'b0000;
    GSharePlugin_logic_mem_counter[6754] = 4'b0000;
    GSharePlugin_logic_mem_counter[6755] = 4'b0000;
    GSharePlugin_logic_mem_counter[6756] = 4'b0000;
    GSharePlugin_logic_mem_counter[6757] = 4'b0000;
    GSharePlugin_logic_mem_counter[6758] = 4'b0000;
    GSharePlugin_logic_mem_counter[6759] = 4'b0000;
    GSharePlugin_logic_mem_counter[6760] = 4'b0000;
    GSharePlugin_logic_mem_counter[6761] = 4'b0000;
    GSharePlugin_logic_mem_counter[6762] = 4'b0000;
    GSharePlugin_logic_mem_counter[6763] = 4'b0000;
    GSharePlugin_logic_mem_counter[6764] = 4'b0000;
    GSharePlugin_logic_mem_counter[6765] = 4'b0000;
    GSharePlugin_logic_mem_counter[6766] = 4'b0000;
    GSharePlugin_logic_mem_counter[6767] = 4'b0000;
    GSharePlugin_logic_mem_counter[6768] = 4'b0000;
    GSharePlugin_logic_mem_counter[6769] = 4'b0000;
    GSharePlugin_logic_mem_counter[6770] = 4'b0000;
    GSharePlugin_logic_mem_counter[6771] = 4'b0000;
    GSharePlugin_logic_mem_counter[6772] = 4'b0000;
    GSharePlugin_logic_mem_counter[6773] = 4'b0000;
    GSharePlugin_logic_mem_counter[6774] = 4'b0000;
    GSharePlugin_logic_mem_counter[6775] = 4'b0000;
    GSharePlugin_logic_mem_counter[6776] = 4'b0000;
    GSharePlugin_logic_mem_counter[6777] = 4'b0000;
    GSharePlugin_logic_mem_counter[6778] = 4'b0000;
    GSharePlugin_logic_mem_counter[6779] = 4'b0000;
    GSharePlugin_logic_mem_counter[6780] = 4'b0000;
    GSharePlugin_logic_mem_counter[6781] = 4'b0000;
    GSharePlugin_logic_mem_counter[6782] = 4'b0000;
    GSharePlugin_logic_mem_counter[6783] = 4'b0000;
    GSharePlugin_logic_mem_counter[6784] = 4'b0000;
    GSharePlugin_logic_mem_counter[6785] = 4'b0000;
    GSharePlugin_logic_mem_counter[6786] = 4'b0000;
    GSharePlugin_logic_mem_counter[6787] = 4'b0000;
    GSharePlugin_logic_mem_counter[6788] = 4'b0000;
    GSharePlugin_logic_mem_counter[6789] = 4'b0000;
    GSharePlugin_logic_mem_counter[6790] = 4'b0000;
    GSharePlugin_logic_mem_counter[6791] = 4'b0000;
    GSharePlugin_logic_mem_counter[6792] = 4'b0000;
    GSharePlugin_logic_mem_counter[6793] = 4'b0000;
    GSharePlugin_logic_mem_counter[6794] = 4'b0000;
    GSharePlugin_logic_mem_counter[6795] = 4'b0000;
    GSharePlugin_logic_mem_counter[6796] = 4'b0000;
    GSharePlugin_logic_mem_counter[6797] = 4'b0000;
    GSharePlugin_logic_mem_counter[6798] = 4'b0000;
    GSharePlugin_logic_mem_counter[6799] = 4'b0000;
    GSharePlugin_logic_mem_counter[6800] = 4'b0000;
    GSharePlugin_logic_mem_counter[6801] = 4'b0000;
    GSharePlugin_logic_mem_counter[6802] = 4'b0000;
    GSharePlugin_logic_mem_counter[6803] = 4'b0000;
    GSharePlugin_logic_mem_counter[6804] = 4'b0000;
    GSharePlugin_logic_mem_counter[6805] = 4'b0000;
    GSharePlugin_logic_mem_counter[6806] = 4'b0000;
    GSharePlugin_logic_mem_counter[6807] = 4'b0000;
    GSharePlugin_logic_mem_counter[6808] = 4'b0000;
    GSharePlugin_logic_mem_counter[6809] = 4'b0000;
    GSharePlugin_logic_mem_counter[6810] = 4'b0000;
    GSharePlugin_logic_mem_counter[6811] = 4'b0000;
    GSharePlugin_logic_mem_counter[6812] = 4'b0000;
    GSharePlugin_logic_mem_counter[6813] = 4'b0000;
    GSharePlugin_logic_mem_counter[6814] = 4'b0000;
    GSharePlugin_logic_mem_counter[6815] = 4'b0000;
    GSharePlugin_logic_mem_counter[6816] = 4'b0000;
    GSharePlugin_logic_mem_counter[6817] = 4'b0000;
    GSharePlugin_logic_mem_counter[6818] = 4'b0000;
    GSharePlugin_logic_mem_counter[6819] = 4'b0000;
    GSharePlugin_logic_mem_counter[6820] = 4'b0000;
    GSharePlugin_logic_mem_counter[6821] = 4'b0000;
    GSharePlugin_logic_mem_counter[6822] = 4'b0000;
    GSharePlugin_logic_mem_counter[6823] = 4'b0000;
    GSharePlugin_logic_mem_counter[6824] = 4'b0000;
    GSharePlugin_logic_mem_counter[6825] = 4'b0000;
    GSharePlugin_logic_mem_counter[6826] = 4'b0000;
    GSharePlugin_logic_mem_counter[6827] = 4'b0000;
    GSharePlugin_logic_mem_counter[6828] = 4'b0000;
    GSharePlugin_logic_mem_counter[6829] = 4'b0000;
    GSharePlugin_logic_mem_counter[6830] = 4'b0000;
    GSharePlugin_logic_mem_counter[6831] = 4'b0000;
    GSharePlugin_logic_mem_counter[6832] = 4'b0000;
    GSharePlugin_logic_mem_counter[6833] = 4'b0000;
    GSharePlugin_logic_mem_counter[6834] = 4'b0000;
    GSharePlugin_logic_mem_counter[6835] = 4'b0000;
    GSharePlugin_logic_mem_counter[6836] = 4'b0000;
    GSharePlugin_logic_mem_counter[6837] = 4'b0000;
    GSharePlugin_logic_mem_counter[6838] = 4'b0000;
    GSharePlugin_logic_mem_counter[6839] = 4'b0000;
    GSharePlugin_logic_mem_counter[6840] = 4'b0000;
    GSharePlugin_logic_mem_counter[6841] = 4'b0000;
    GSharePlugin_logic_mem_counter[6842] = 4'b0000;
    GSharePlugin_logic_mem_counter[6843] = 4'b0000;
    GSharePlugin_logic_mem_counter[6844] = 4'b0000;
    GSharePlugin_logic_mem_counter[6845] = 4'b0000;
    GSharePlugin_logic_mem_counter[6846] = 4'b0000;
    GSharePlugin_logic_mem_counter[6847] = 4'b0000;
    GSharePlugin_logic_mem_counter[6848] = 4'b0000;
    GSharePlugin_logic_mem_counter[6849] = 4'b0000;
    GSharePlugin_logic_mem_counter[6850] = 4'b0000;
    GSharePlugin_logic_mem_counter[6851] = 4'b0000;
    GSharePlugin_logic_mem_counter[6852] = 4'b0000;
    GSharePlugin_logic_mem_counter[6853] = 4'b0000;
    GSharePlugin_logic_mem_counter[6854] = 4'b0000;
    GSharePlugin_logic_mem_counter[6855] = 4'b0000;
    GSharePlugin_logic_mem_counter[6856] = 4'b0000;
    GSharePlugin_logic_mem_counter[6857] = 4'b0000;
    GSharePlugin_logic_mem_counter[6858] = 4'b0000;
    GSharePlugin_logic_mem_counter[6859] = 4'b0000;
    GSharePlugin_logic_mem_counter[6860] = 4'b0000;
    GSharePlugin_logic_mem_counter[6861] = 4'b0000;
    GSharePlugin_logic_mem_counter[6862] = 4'b0000;
    GSharePlugin_logic_mem_counter[6863] = 4'b0000;
    GSharePlugin_logic_mem_counter[6864] = 4'b0000;
    GSharePlugin_logic_mem_counter[6865] = 4'b0000;
    GSharePlugin_logic_mem_counter[6866] = 4'b0000;
    GSharePlugin_logic_mem_counter[6867] = 4'b0000;
    GSharePlugin_logic_mem_counter[6868] = 4'b0000;
    GSharePlugin_logic_mem_counter[6869] = 4'b0000;
    GSharePlugin_logic_mem_counter[6870] = 4'b0000;
    GSharePlugin_logic_mem_counter[6871] = 4'b0000;
    GSharePlugin_logic_mem_counter[6872] = 4'b0000;
    GSharePlugin_logic_mem_counter[6873] = 4'b0000;
    GSharePlugin_logic_mem_counter[6874] = 4'b0000;
    GSharePlugin_logic_mem_counter[6875] = 4'b0000;
    GSharePlugin_logic_mem_counter[6876] = 4'b0000;
    GSharePlugin_logic_mem_counter[6877] = 4'b0000;
    GSharePlugin_logic_mem_counter[6878] = 4'b0000;
    GSharePlugin_logic_mem_counter[6879] = 4'b0000;
    GSharePlugin_logic_mem_counter[6880] = 4'b0000;
    GSharePlugin_logic_mem_counter[6881] = 4'b0000;
    GSharePlugin_logic_mem_counter[6882] = 4'b0000;
    GSharePlugin_logic_mem_counter[6883] = 4'b0000;
    GSharePlugin_logic_mem_counter[6884] = 4'b0000;
    GSharePlugin_logic_mem_counter[6885] = 4'b0000;
    GSharePlugin_logic_mem_counter[6886] = 4'b0000;
    GSharePlugin_logic_mem_counter[6887] = 4'b0000;
    GSharePlugin_logic_mem_counter[6888] = 4'b0000;
    GSharePlugin_logic_mem_counter[6889] = 4'b0000;
    GSharePlugin_logic_mem_counter[6890] = 4'b0000;
    GSharePlugin_logic_mem_counter[6891] = 4'b0000;
    GSharePlugin_logic_mem_counter[6892] = 4'b0000;
    GSharePlugin_logic_mem_counter[6893] = 4'b0000;
    GSharePlugin_logic_mem_counter[6894] = 4'b0000;
    GSharePlugin_logic_mem_counter[6895] = 4'b0000;
    GSharePlugin_logic_mem_counter[6896] = 4'b0000;
    GSharePlugin_logic_mem_counter[6897] = 4'b0000;
    GSharePlugin_logic_mem_counter[6898] = 4'b0000;
    GSharePlugin_logic_mem_counter[6899] = 4'b0000;
    GSharePlugin_logic_mem_counter[6900] = 4'b0000;
    GSharePlugin_logic_mem_counter[6901] = 4'b0000;
    GSharePlugin_logic_mem_counter[6902] = 4'b0000;
    GSharePlugin_logic_mem_counter[6903] = 4'b0000;
    GSharePlugin_logic_mem_counter[6904] = 4'b0000;
    GSharePlugin_logic_mem_counter[6905] = 4'b0000;
    GSharePlugin_logic_mem_counter[6906] = 4'b0000;
    GSharePlugin_logic_mem_counter[6907] = 4'b0000;
    GSharePlugin_logic_mem_counter[6908] = 4'b0000;
    GSharePlugin_logic_mem_counter[6909] = 4'b0000;
    GSharePlugin_logic_mem_counter[6910] = 4'b0000;
    GSharePlugin_logic_mem_counter[6911] = 4'b0000;
    GSharePlugin_logic_mem_counter[6912] = 4'b0000;
    GSharePlugin_logic_mem_counter[6913] = 4'b0000;
    GSharePlugin_logic_mem_counter[6914] = 4'b0000;
    GSharePlugin_logic_mem_counter[6915] = 4'b0000;
    GSharePlugin_logic_mem_counter[6916] = 4'b0000;
    GSharePlugin_logic_mem_counter[6917] = 4'b0000;
    GSharePlugin_logic_mem_counter[6918] = 4'b0000;
    GSharePlugin_logic_mem_counter[6919] = 4'b0000;
    GSharePlugin_logic_mem_counter[6920] = 4'b0000;
    GSharePlugin_logic_mem_counter[6921] = 4'b0000;
    GSharePlugin_logic_mem_counter[6922] = 4'b0000;
    GSharePlugin_logic_mem_counter[6923] = 4'b0000;
    GSharePlugin_logic_mem_counter[6924] = 4'b0000;
    GSharePlugin_logic_mem_counter[6925] = 4'b0000;
    GSharePlugin_logic_mem_counter[6926] = 4'b0000;
    GSharePlugin_logic_mem_counter[6927] = 4'b0000;
    GSharePlugin_logic_mem_counter[6928] = 4'b0000;
    GSharePlugin_logic_mem_counter[6929] = 4'b0000;
    GSharePlugin_logic_mem_counter[6930] = 4'b0000;
    GSharePlugin_logic_mem_counter[6931] = 4'b0000;
    GSharePlugin_logic_mem_counter[6932] = 4'b0000;
    GSharePlugin_logic_mem_counter[6933] = 4'b0000;
    GSharePlugin_logic_mem_counter[6934] = 4'b0000;
    GSharePlugin_logic_mem_counter[6935] = 4'b0000;
    GSharePlugin_logic_mem_counter[6936] = 4'b0000;
    GSharePlugin_logic_mem_counter[6937] = 4'b0000;
    GSharePlugin_logic_mem_counter[6938] = 4'b0000;
    GSharePlugin_logic_mem_counter[6939] = 4'b0000;
    GSharePlugin_logic_mem_counter[6940] = 4'b0000;
    GSharePlugin_logic_mem_counter[6941] = 4'b0000;
    GSharePlugin_logic_mem_counter[6942] = 4'b0000;
    GSharePlugin_logic_mem_counter[6943] = 4'b0000;
    GSharePlugin_logic_mem_counter[6944] = 4'b0000;
    GSharePlugin_logic_mem_counter[6945] = 4'b0000;
    GSharePlugin_logic_mem_counter[6946] = 4'b0000;
    GSharePlugin_logic_mem_counter[6947] = 4'b0000;
    GSharePlugin_logic_mem_counter[6948] = 4'b0000;
    GSharePlugin_logic_mem_counter[6949] = 4'b0000;
    GSharePlugin_logic_mem_counter[6950] = 4'b0000;
    GSharePlugin_logic_mem_counter[6951] = 4'b0000;
    GSharePlugin_logic_mem_counter[6952] = 4'b0000;
    GSharePlugin_logic_mem_counter[6953] = 4'b0000;
    GSharePlugin_logic_mem_counter[6954] = 4'b0000;
    GSharePlugin_logic_mem_counter[6955] = 4'b0000;
    GSharePlugin_logic_mem_counter[6956] = 4'b0000;
    GSharePlugin_logic_mem_counter[6957] = 4'b0000;
    GSharePlugin_logic_mem_counter[6958] = 4'b0000;
    GSharePlugin_logic_mem_counter[6959] = 4'b0000;
    GSharePlugin_logic_mem_counter[6960] = 4'b0000;
    GSharePlugin_logic_mem_counter[6961] = 4'b0000;
    GSharePlugin_logic_mem_counter[6962] = 4'b0000;
    GSharePlugin_logic_mem_counter[6963] = 4'b0000;
    GSharePlugin_logic_mem_counter[6964] = 4'b0000;
    GSharePlugin_logic_mem_counter[6965] = 4'b0000;
    GSharePlugin_logic_mem_counter[6966] = 4'b0000;
    GSharePlugin_logic_mem_counter[6967] = 4'b0000;
    GSharePlugin_logic_mem_counter[6968] = 4'b0000;
    GSharePlugin_logic_mem_counter[6969] = 4'b0000;
    GSharePlugin_logic_mem_counter[6970] = 4'b0000;
    GSharePlugin_logic_mem_counter[6971] = 4'b0000;
    GSharePlugin_logic_mem_counter[6972] = 4'b0000;
    GSharePlugin_logic_mem_counter[6973] = 4'b0000;
    GSharePlugin_logic_mem_counter[6974] = 4'b0000;
    GSharePlugin_logic_mem_counter[6975] = 4'b0000;
    GSharePlugin_logic_mem_counter[6976] = 4'b0000;
    GSharePlugin_logic_mem_counter[6977] = 4'b0000;
    GSharePlugin_logic_mem_counter[6978] = 4'b0000;
    GSharePlugin_logic_mem_counter[6979] = 4'b0000;
    GSharePlugin_logic_mem_counter[6980] = 4'b0000;
    GSharePlugin_logic_mem_counter[6981] = 4'b0000;
    GSharePlugin_logic_mem_counter[6982] = 4'b0000;
    GSharePlugin_logic_mem_counter[6983] = 4'b0000;
    GSharePlugin_logic_mem_counter[6984] = 4'b0000;
    GSharePlugin_logic_mem_counter[6985] = 4'b0000;
    GSharePlugin_logic_mem_counter[6986] = 4'b0000;
    GSharePlugin_logic_mem_counter[6987] = 4'b0000;
    GSharePlugin_logic_mem_counter[6988] = 4'b0000;
    GSharePlugin_logic_mem_counter[6989] = 4'b0000;
    GSharePlugin_logic_mem_counter[6990] = 4'b0000;
    GSharePlugin_logic_mem_counter[6991] = 4'b0000;
    GSharePlugin_logic_mem_counter[6992] = 4'b0000;
    GSharePlugin_logic_mem_counter[6993] = 4'b0000;
    GSharePlugin_logic_mem_counter[6994] = 4'b0000;
    GSharePlugin_logic_mem_counter[6995] = 4'b0000;
    GSharePlugin_logic_mem_counter[6996] = 4'b0000;
    GSharePlugin_logic_mem_counter[6997] = 4'b0000;
    GSharePlugin_logic_mem_counter[6998] = 4'b0000;
    GSharePlugin_logic_mem_counter[6999] = 4'b0000;
    GSharePlugin_logic_mem_counter[7000] = 4'b0000;
    GSharePlugin_logic_mem_counter[7001] = 4'b0000;
    GSharePlugin_logic_mem_counter[7002] = 4'b0000;
    GSharePlugin_logic_mem_counter[7003] = 4'b0000;
    GSharePlugin_logic_mem_counter[7004] = 4'b0000;
    GSharePlugin_logic_mem_counter[7005] = 4'b0000;
    GSharePlugin_logic_mem_counter[7006] = 4'b0000;
    GSharePlugin_logic_mem_counter[7007] = 4'b0000;
    GSharePlugin_logic_mem_counter[7008] = 4'b0000;
    GSharePlugin_logic_mem_counter[7009] = 4'b0000;
    GSharePlugin_logic_mem_counter[7010] = 4'b0000;
    GSharePlugin_logic_mem_counter[7011] = 4'b0000;
    GSharePlugin_logic_mem_counter[7012] = 4'b0000;
    GSharePlugin_logic_mem_counter[7013] = 4'b0000;
    GSharePlugin_logic_mem_counter[7014] = 4'b0000;
    GSharePlugin_logic_mem_counter[7015] = 4'b0000;
    GSharePlugin_logic_mem_counter[7016] = 4'b0000;
    GSharePlugin_logic_mem_counter[7017] = 4'b0000;
    GSharePlugin_logic_mem_counter[7018] = 4'b0000;
    GSharePlugin_logic_mem_counter[7019] = 4'b0000;
    GSharePlugin_logic_mem_counter[7020] = 4'b0000;
    GSharePlugin_logic_mem_counter[7021] = 4'b0000;
    GSharePlugin_logic_mem_counter[7022] = 4'b0000;
    GSharePlugin_logic_mem_counter[7023] = 4'b0000;
    GSharePlugin_logic_mem_counter[7024] = 4'b0000;
    GSharePlugin_logic_mem_counter[7025] = 4'b0000;
    GSharePlugin_logic_mem_counter[7026] = 4'b0000;
    GSharePlugin_logic_mem_counter[7027] = 4'b0000;
    GSharePlugin_logic_mem_counter[7028] = 4'b0000;
    GSharePlugin_logic_mem_counter[7029] = 4'b0000;
    GSharePlugin_logic_mem_counter[7030] = 4'b0000;
    GSharePlugin_logic_mem_counter[7031] = 4'b0000;
    GSharePlugin_logic_mem_counter[7032] = 4'b0000;
    GSharePlugin_logic_mem_counter[7033] = 4'b0000;
    GSharePlugin_logic_mem_counter[7034] = 4'b0000;
    GSharePlugin_logic_mem_counter[7035] = 4'b0000;
    GSharePlugin_logic_mem_counter[7036] = 4'b0000;
    GSharePlugin_logic_mem_counter[7037] = 4'b0000;
    GSharePlugin_logic_mem_counter[7038] = 4'b0000;
    GSharePlugin_logic_mem_counter[7039] = 4'b0000;
    GSharePlugin_logic_mem_counter[7040] = 4'b0000;
    GSharePlugin_logic_mem_counter[7041] = 4'b0000;
    GSharePlugin_logic_mem_counter[7042] = 4'b0000;
    GSharePlugin_logic_mem_counter[7043] = 4'b0000;
    GSharePlugin_logic_mem_counter[7044] = 4'b0000;
    GSharePlugin_logic_mem_counter[7045] = 4'b0000;
    GSharePlugin_logic_mem_counter[7046] = 4'b0000;
    GSharePlugin_logic_mem_counter[7047] = 4'b0000;
    GSharePlugin_logic_mem_counter[7048] = 4'b0000;
    GSharePlugin_logic_mem_counter[7049] = 4'b0000;
    GSharePlugin_logic_mem_counter[7050] = 4'b0000;
    GSharePlugin_logic_mem_counter[7051] = 4'b0000;
    GSharePlugin_logic_mem_counter[7052] = 4'b0000;
    GSharePlugin_logic_mem_counter[7053] = 4'b0000;
    GSharePlugin_logic_mem_counter[7054] = 4'b0000;
    GSharePlugin_logic_mem_counter[7055] = 4'b0000;
    GSharePlugin_logic_mem_counter[7056] = 4'b0000;
    GSharePlugin_logic_mem_counter[7057] = 4'b0000;
    GSharePlugin_logic_mem_counter[7058] = 4'b0000;
    GSharePlugin_logic_mem_counter[7059] = 4'b0000;
    GSharePlugin_logic_mem_counter[7060] = 4'b0000;
    GSharePlugin_logic_mem_counter[7061] = 4'b0000;
    GSharePlugin_logic_mem_counter[7062] = 4'b0000;
    GSharePlugin_logic_mem_counter[7063] = 4'b0000;
    GSharePlugin_logic_mem_counter[7064] = 4'b0000;
    GSharePlugin_logic_mem_counter[7065] = 4'b0000;
    GSharePlugin_logic_mem_counter[7066] = 4'b0000;
    GSharePlugin_logic_mem_counter[7067] = 4'b0000;
    GSharePlugin_logic_mem_counter[7068] = 4'b0000;
    GSharePlugin_logic_mem_counter[7069] = 4'b0000;
    GSharePlugin_logic_mem_counter[7070] = 4'b0000;
    GSharePlugin_logic_mem_counter[7071] = 4'b0000;
    GSharePlugin_logic_mem_counter[7072] = 4'b0000;
    GSharePlugin_logic_mem_counter[7073] = 4'b0000;
    GSharePlugin_logic_mem_counter[7074] = 4'b0000;
    GSharePlugin_logic_mem_counter[7075] = 4'b0000;
    GSharePlugin_logic_mem_counter[7076] = 4'b0000;
    GSharePlugin_logic_mem_counter[7077] = 4'b0000;
    GSharePlugin_logic_mem_counter[7078] = 4'b0000;
    GSharePlugin_logic_mem_counter[7079] = 4'b0000;
    GSharePlugin_logic_mem_counter[7080] = 4'b0000;
    GSharePlugin_logic_mem_counter[7081] = 4'b0000;
    GSharePlugin_logic_mem_counter[7082] = 4'b0000;
    GSharePlugin_logic_mem_counter[7083] = 4'b0000;
    GSharePlugin_logic_mem_counter[7084] = 4'b0000;
    GSharePlugin_logic_mem_counter[7085] = 4'b0000;
    GSharePlugin_logic_mem_counter[7086] = 4'b0000;
    GSharePlugin_logic_mem_counter[7087] = 4'b0000;
    GSharePlugin_logic_mem_counter[7088] = 4'b0000;
    GSharePlugin_logic_mem_counter[7089] = 4'b0000;
    GSharePlugin_logic_mem_counter[7090] = 4'b0000;
    GSharePlugin_logic_mem_counter[7091] = 4'b0000;
    GSharePlugin_logic_mem_counter[7092] = 4'b0000;
    GSharePlugin_logic_mem_counter[7093] = 4'b0000;
    GSharePlugin_logic_mem_counter[7094] = 4'b0000;
    GSharePlugin_logic_mem_counter[7095] = 4'b0000;
    GSharePlugin_logic_mem_counter[7096] = 4'b0000;
    GSharePlugin_logic_mem_counter[7097] = 4'b0000;
    GSharePlugin_logic_mem_counter[7098] = 4'b0000;
    GSharePlugin_logic_mem_counter[7099] = 4'b0000;
    GSharePlugin_logic_mem_counter[7100] = 4'b0000;
    GSharePlugin_logic_mem_counter[7101] = 4'b0000;
    GSharePlugin_logic_mem_counter[7102] = 4'b0000;
    GSharePlugin_logic_mem_counter[7103] = 4'b0000;
    GSharePlugin_logic_mem_counter[7104] = 4'b0000;
    GSharePlugin_logic_mem_counter[7105] = 4'b0000;
    GSharePlugin_logic_mem_counter[7106] = 4'b0000;
    GSharePlugin_logic_mem_counter[7107] = 4'b0000;
    GSharePlugin_logic_mem_counter[7108] = 4'b0000;
    GSharePlugin_logic_mem_counter[7109] = 4'b0000;
    GSharePlugin_logic_mem_counter[7110] = 4'b0000;
    GSharePlugin_logic_mem_counter[7111] = 4'b0000;
    GSharePlugin_logic_mem_counter[7112] = 4'b0000;
    GSharePlugin_logic_mem_counter[7113] = 4'b0000;
    GSharePlugin_logic_mem_counter[7114] = 4'b0000;
    GSharePlugin_logic_mem_counter[7115] = 4'b0000;
    GSharePlugin_logic_mem_counter[7116] = 4'b0000;
    GSharePlugin_logic_mem_counter[7117] = 4'b0000;
    GSharePlugin_logic_mem_counter[7118] = 4'b0000;
    GSharePlugin_logic_mem_counter[7119] = 4'b0000;
    GSharePlugin_logic_mem_counter[7120] = 4'b0000;
    GSharePlugin_logic_mem_counter[7121] = 4'b0000;
    GSharePlugin_logic_mem_counter[7122] = 4'b0000;
    GSharePlugin_logic_mem_counter[7123] = 4'b0000;
    GSharePlugin_logic_mem_counter[7124] = 4'b0000;
    GSharePlugin_logic_mem_counter[7125] = 4'b0000;
    GSharePlugin_logic_mem_counter[7126] = 4'b0000;
    GSharePlugin_logic_mem_counter[7127] = 4'b0000;
    GSharePlugin_logic_mem_counter[7128] = 4'b0000;
    GSharePlugin_logic_mem_counter[7129] = 4'b0000;
    GSharePlugin_logic_mem_counter[7130] = 4'b0000;
    GSharePlugin_logic_mem_counter[7131] = 4'b0000;
    GSharePlugin_logic_mem_counter[7132] = 4'b0000;
    GSharePlugin_logic_mem_counter[7133] = 4'b0000;
    GSharePlugin_logic_mem_counter[7134] = 4'b0000;
    GSharePlugin_logic_mem_counter[7135] = 4'b0000;
    GSharePlugin_logic_mem_counter[7136] = 4'b0000;
    GSharePlugin_logic_mem_counter[7137] = 4'b0000;
    GSharePlugin_logic_mem_counter[7138] = 4'b0000;
    GSharePlugin_logic_mem_counter[7139] = 4'b0000;
    GSharePlugin_logic_mem_counter[7140] = 4'b0000;
    GSharePlugin_logic_mem_counter[7141] = 4'b0000;
    GSharePlugin_logic_mem_counter[7142] = 4'b0000;
    GSharePlugin_logic_mem_counter[7143] = 4'b0000;
    GSharePlugin_logic_mem_counter[7144] = 4'b0000;
    GSharePlugin_logic_mem_counter[7145] = 4'b0000;
    GSharePlugin_logic_mem_counter[7146] = 4'b0000;
    GSharePlugin_logic_mem_counter[7147] = 4'b0000;
    GSharePlugin_logic_mem_counter[7148] = 4'b0000;
    GSharePlugin_logic_mem_counter[7149] = 4'b0000;
    GSharePlugin_logic_mem_counter[7150] = 4'b0000;
    GSharePlugin_logic_mem_counter[7151] = 4'b0000;
    GSharePlugin_logic_mem_counter[7152] = 4'b0000;
    GSharePlugin_logic_mem_counter[7153] = 4'b0000;
    GSharePlugin_logic_mem_counter[7154] = 4'b0000;
    GSharePlugin_logic_mem_counter[7155] = 4'b0000;
    GSharePlugin_logic_mem_counter[7156] = 4'b0000;
    GSharePlugin_logic_mem_counter[7157] = 4'b0000;
    GSharePlugin_logic_mem_counter[7158] = 4'b0000;
    GSharePlugin_logic_mem_counter[7159] = 4'b0000;
    GSharePlugin_logic_mem_counter[7160] = 4'b0000;
    GSharePlugin_logic_mem_counter[7161] = 4'b0000;
    GSharePlugin_logic_mem_counter[7162] = 4'b0000;
    GSharePlugin_logic_mem_counter[7163] = 4'b0000;
    GSharePlugin_logic_mem_counter[7164] = 4'b0000;
    GSharePlugin_logic_mem_counter[7165] = 4'b0000;
    GSharePlugin_logic_mem_counter[7166] = 4'b0000;
    GSharePlugin_logic_mem_counter[7167] = 4'b0000;
    GSharePlugin_logic_mem_counter[7168] = 4'b0000;
    GSharePlugin_logic_mem_counter[7169] = 4'b0000;
    GSharePlugin_logic_mem_counter[7170] = 4'b0000;
    GSharePlugin_logic_mem_counter[7171] = 4'b0000;
    GSharePlugin_logic_mem_counter[7172] = 4'b0000;
    GSharePlugin_logic_mem_counter[7173] = 4'b0000;
    GSharePlugin_logic_mem_counter[7174] = 4'b0000;
    GSharePlugin_logic_mem_counter[7175] = 4'b0000;
    GSharePlugin_logic_mem_counter[7176] = 4'b0000;
    GSharePlugin_logic_mem_counter[7177] = 4'b0000;
    GSharePlugin_logic_mem_counter[7178] = 4'b0000;
    GSharePlugin_logic_mem_counter[7179] = 4'b0000;
    GSharePlugin_logic_mem_counter[7180] = 4'b0000;
    GSharePlugin_logic_mem_counter[7181] = 4'b0000;
    GSharePlugin_logic_mem_counter[7182] = 4'b0000;
    GSharePlugin_logic_mem_counter[7183] = 4'b0000;
    GSharePlugin_logic_mem_counter[7184] = 4'b0000;
    GSharePlugin_logic_mem_counter[7185] = 4'b0000;
    GSharePlugin_logic_mem_counter[7186] = 4'b0000;
    GSharePlugin_logic_mem_counter[7187] = 4'b0000;
    GSharePlugin_logic_mem_counter[7188] = 4'b0000;
    GSharePlugin_logic_mem_counter[7189] = 4'b0000;
    GSharePlugin_logic_mem_counter[7190] = 4'b0000;
    GSharePlugin_logic_mem_counter[7191] = 4'b0000;
    GSharePlugin_logic_mem_counter[7192] = 4'b0000;
    GSharePlugin_logic_mem_counter[7193] = 4'b0000;
    GSharePlugin_logic_mem_counter[7194] = 4'b0000;
    GSharePlugin_logic_mem_counter[7195] = 4'b0000;
    GSharePlugin_logic_mem_counter[7196] = 4'b0000;
    GSharePlugin_logic_mem_counter[7197] = 4'b0000;
    GSharePlugin_logic_mem_counter[7198] = 4'b0000;
    GSharePlugin_logic_mem_counter[7199] = 4'b0000;
    GSharePlugin_logic_mem_counter[7200] = 4'b0000;
    GSharePlugin_logic_mem_counter[7201] = 4'b0000;
    GSharePlugin_logic_mem_counter[7202] = 4'b0000;
    GSharePlugin_logic_mem_counter[7203] = 4'b0000;
    GSharePlugin_logic_mem_counter[7204] = 4'b0000;
    GSharePlugin_logic_mem_counter[7205] = 4'b0000;
    GSharePlugin_logic_mem_counter[7206] = 4'b0000;
    GSharePlugin_logic_mem_counter[7207] = 4'b0000;
    GSharePlugin_logic_mem_counter[7208] = 4'b0000;
    GSharePlugin_logic_mem_counter[7209] = 4'b0000;
    GSharePlugin_logic_mem_counter[7210] = 4'b0000;
    GSharePlugin_logic_mem_counter[7211] = 4'b0000;
    GSharePlugin_logic_mem_counter[7212] = 4'b0000;
    GSharePlugin_logic_mem_counter[7213] = 4'b0000;
    GSharePlugin_logic_mem_counter[7214] = 4'b0000;
    GSharePlugin_logic_mem_counter[7215] = 4'b0000;
    GSharePlugin_logic_mem_counter[7216] = 4'b0000;
    GSharePlugin_logic_mem_counter[7217] = 4'b0000;
    GSharePlugin_logic_mem_counter[7218] = 4'b0000;
    GSharePlugin_logic_mem_counter[7219] = 4'b0000;
    GSharePlugin_logic_mem_counter[7220] = 4'b0000;
    GSharePlugin_logic_mem_counter[7221] = 4'b0000;
    GSharePlugin_logic_mem_counter[7222] = 4'b0000;
    GSharePlugin_logic_mem_counter[7223] = 4'b0000;
    GSharePlugin_logic_mem_counter[7224] = 4'b0000;
    GSharePlugin_logic_mem_counter[7225] = 4'b0000;
    GSharePlugin_logic_mem_counter[7226] = 4'b0000;
    GSharePlugin_logic_mem_counter[7227] = 4'b0000;
    GSharePlugin_logic_mem_counter[7228] = 4'b0000;
    GSharePlugin_logic_mem_counter[7229] = 4'b0000;
    GSharePlugin_logic_mem_counter[7230] = 4'b0000;
    GSharePlugin_logic_mem_counter[7231] = 4'b0000;
    GSharePlugin_logic_mem_counter[7232] = 4'b0000;
    GSharePlugin_logic_mem_counter[7233] = 4'b0000;
    GSharePlugin_logic_mem_counter[7234] = 4'b0000;
    GSharePlugin_logic_mem_counter[7235] = 4'b0000;
    GSharePlugin_logic_mem_counter[7236] = 4'b0000;
    GSharePlugin_logic_mem_counter[7237] = 4'b0000;
    GSharePlugin_logic_mem_counter[7238] = 4'b0000;
    GSharePlugin_logic_mem_counter[7239] = 4'b0000;
    GSharePlugin_logic_mem_counter[7240] = 4'b0000;
    GSharePlugin_logic_mem_counter[7241] = 4'b0000;
    GSharePlugin_logic_mem_counter[7242] = 4'b0000;
    GSharePlugin_logic_mem_counter[7243] = 4'b0000;
    GSharePlugin_logic_mem_counter[7244] = 4'b0000;
    GSharePlugin_logic_mem_counter[7245] = 4'b0000;
    GSharePlugin_logic_mem_counter[7246] = 4'b0000;
    GSharePlugin_logic_mem_counter[7247] = 4'b0000;
    GSharePlugin_logic_mem_counter[7248] = 4'b0000;
    GSharePlugin_logic_mem_counter[7249] = 4'b0000;
    GSharePlugin_logic_mem_counter[7250] = 4'b0000;
    GSharePlugin_logic_mem_counter[7251] = 4'b0000;
    GSharePlugin_logic_mem_counter[7252] = 4'b0000;
    GSharePlugin_logic_mem_counter[7253] = 4'b0000;
    GSharePlugin_logic_mem_counter[7254] = 4'b0000;
    GSharePlugin_logic_mem_counter[7255] = 4'b0000;
    GSharePlugin_logic_mem_counter[7256] = 4'b0000;
    GSharePlugin_logic_mem_counter[7257] = 4'b0000;
    GSharePlugin_logic_mem_counter[7258] = 4'b0000;
    GSharePlugin_logic_mem_counter[7259] = 4'b0000;
    GSharePlugin_logic_mem_counter[7260] = 4'b0000;
    GSharePlugin_logic_mem_counter[7261] = 4'b0000;
    GSharePlugin_logic_mem_counter[7262] = 4'b0000;
    GSharePlugin_logic_mem_counter[7263] = 4'b0000;
    GSharePlugin_logic_mem_counter[7264] = 4'b0000;
    GSharePlugin_logic_mem_counter[7265] = 4'b0000;
    GSharePlugin_logic_mem_counter[7266] = 4'b0000;
    GSharePlugin_logic_mem_counter[7267] = 4'b0000;
    GSharePlugin_logic_mem_counter[7268] = 4'b0000;
    GSharePlugin_logic_mem_counter[7269] = 4'b0000;
    GSharePlugin_logic_mem_counter[7270] = 4'b0000;
    GSharePlugin_logic_mem_counter[7271] = 4'b0000;
    GSharePlugin_logic_mem_counter[7272] = 4'b0000;
    GSharePlugin_logic_mem_counter[7273] = 4'b0000;
    GSharePlugin_logic_mem_counter[7274] = 4'b0000;
    GSharePlugin_logic_mem_counter[7275] = 4'b0000;
    GSharePlugin_logic_mem_counter[7276] = 4'b0000;
    GSharePlugin_logic_mem_counter[7277] = 4'b0000;
    GSharePlugin_logic_mem_counter[7278] = 4'b0000;
    GSharePlugin_logic_mem_counter[7279] = 4'b0000;
    GSharePlugin_logic_mem_counter[7280] = 4'b0000;
    GSharePlugin_logic_mem_counter[7281] = 4'b0000;
    GSharePlugin_logic_mem_counter[7282] = 4'b0000;
    GSharePlugin_logic_mem_counter[7283] = 4'b0000;
    GSharePlugin_logic_mem_counter[7284] = 4'b0000;
    GSharePlugin_logic_mem_counter[7285] = 4'b0000;
    GSharePlugin_logic_mem_counter[7286] = 4'b0000;
    GSharePlugin_logic_mem_counter[7287] = 4'b0000;
    GSharePlugin_logic_mem_counter[7288] = 4'b0000;
    GSharePlugin_logic_mem_counter[7289] = 4'b0000;
    GSharePlugin_logic_mem_counter[7290] = 4'b0000;
    GSharePlugin_logic_mem_counter[7291] = 4'b0000;
    GSharePlugin_logic_mem_counter[7292] = 4'b0000;
    GSharePlugin_logic_mem_counter[7293] = 4'b0000;
    GSharePlugin_logic_mem_counter[7294] = 4'b0000;
    GSharePlugin_logic_mem_counter[7295] = 4'b0000;
    GSharePlugin_logic_mem_counter[7296] = 4'b0000;
    GSharePlugin_logic_mem_counter[7297] = 4'b0000;
    GSharePlugin_logic_mem_counter[7298] = 4'b0000;
    GSharePlugin_logic_mem_counter[7299] = 4'b0000;
    GSharePlugin_logic_mem_counter[7300] = 4'b0000;
    GSharePlugin_logic_mem_counter[7301] = 4'b0000;
    GSharePlugin_logic_mem_counter[7302] = 4'b0000;
    GSharePlugin_logic_mem_counter[7303] = 4'b0000;
    GSharePlugin_logic_mem_counter[7304] = 4'b0000;
    GSharePlugin_logic_mem_counter[7305] = 4'b0000;
    GSharePlugin_logic_mem_counter[7306] = 4'b0000;
    GSharePlugin_logic_mem_counter[7307] = 4'b0000;
    GSharePlugin_logic_mem_counter[7308] = 4'b0000;
    GSharePlugin_logic_mem_counter[7309] = 4'b0000;
    GSharePlugin_logic_mem_counter[7310] = 4'b0000;
    GSharePlugin_logic_mem_counter[7311] = 4'b0000;
    GSharePlugin_logic_mem_counter[7312] = 4'b0000;
    GSharePlugin_logic_mem_counter[7313] = 4'b0000;
    GSharePlugin_logic_mem_counter[7314] = 4'b0000;
    GSharePlugin_logic_mem_counter[7315] = 4'b0000;
    GSharePlugin_logic_mem_counter[7316] = 4'b0000;
    GSharePlugin_logic_mem_counter[7317] = 4'b0000;
    GSharePlugin_logic_mem_counter[7318] = 4'b0000;
    GSharePlugin_logic_mem_counter[7319] = 4'b0000;
    GSharePlugin_logic_mem_counter[7320] = 4'b0000;
    GSharePlugin_logic_mem_counter[7321] = 4'b0000;
    GSharePlugin_logic_mem_counter[7322] = 4'b0000;
    GSharePlugin_logic_mem_counter[7323] = 4'b0000;
    GSharePlugin_logic_mem_counter[7324] = 4'b0000;
    GSharePlugin_logic_mem_counter[7325] = 4'b0000;
    GSharePlugin_logic_mem_counter[7326] = 4'b0000;
    GSharePlugin_logic_mem_counter[7327] = 4'b0000;
    GSharePlugin_logic_mem_counter[7328] = 4'b0000;
    GSharePlugin_logic_mem_counter[7329] = 4'b0000;
    GSharePlugin_logic_mem_counter[7330] = 4'b0000;
    GSharePlugin_logic_mem_counter[7331] = 4'b0000;
    GSharePlugin_logic_mem_counter[7332] = 4'b0000;
    GSharePlugin_logic_mem_counter[7333] = 4'b0000;
    GSharePlugin_logic_mem_counter[7334] = 4'b0000;
    GSharePlugin_logic_mem_counter[7335] = 4'b0000;
    GSharePlugin_logic_mem_counter[7336] = 4'b0000;
    GSharePlugin_logic_mem_counter[7337] = 4'b0000;
    GSharePlugin_logic_mem_counter[7338] = 4'b0000;
    GSharePlugin_logic_mem_counter[7339] = 4'b0000;
    GSharePlugin_logic_mem_counter[7340] = 4'b0000;
    GSharePlugin_logic_mem_counter[7341] = 4'b0000;
    GSharePlugin_logic_mem_counter[7342] = 4'b0000;
    GSharePlugin_logic_mem_counter[7343] = 4'b0000;
    GSharePlugin_logic_mem_counter[7344] = 4'b0000;
    GSharePlugin_logic_mem_counter[7345] = 4'b0000;
    GSharePlugin_logic_mem_counter[7346] = 4'b0000;
    GSharePlugin_logic_mem_counter[7347] = 4'b0000;
    GSharePlugin_logic_mem_counter[7348] = 4'b0000;
    GSharePlugin_logic_mem_counter[7349] = 4'b0000;
    GSharePlugin_logic_mem_counter[7350] = 4'b0000;
    GSharePlugin_logic_mem_counter[7351] = 4'b0000;
    GSharePlugin_logic_mem_counter[7352] = 4'b0000;
    GSharePlugin_logic_mem_counter[7353] = 4'b0000;
    GSharePlugin_logic_mem_counter[7354] = 4'b0000;
    GSharePlugin_logic_mem_counter[7355] = 4'b0000;
    GSharePlugin_logic_mem_counter[7356] = 4'b0000;
    GSharePlugin_logic_mem_counter[7357] = 4'b0000;
    GSharePlugin_logic_mem_counter[7358] = 4'b0000;
    GSharePlugin_logic_mem_counter[7359] = 4'b0000;
    GSharePlugin_logic_mem_counter[7360] = 4'b0000;
    GSharePlugin_logic_mem_counter[7361] = 4'b0000;
    GSharePlugin_logic_mem_counter[7362] = 4'b0000;
    GSharePlugin_logic_mem_counter[7363] = 4'b0000;
    GSharePlugin_logic_mem_counter[7364] = 4'b0000;
    GSharePlugin_logic_mem_counter[7365] = 4'b0000;
    GSharePlugin_logic_mem_counter[7366] = 4'b0000;
    GSharePlugin_logic_mem_counter[7367] = 4'b0000;
    GSharePlugin_logic_mem_counter[7368] = 4'b0000;
    GSharePlugin_logic_mem_counter[7369] = 4'b0000;
    GSharePlugin_logic_mem_counter[7370] = 4'b0000;
    GSharePlugin_logic_mem_counter[7371] = 4'b0000;
    GSharePlugin_logic_mem_counter[7372] = 4'b0000;
    GSharePlugin_logic_mem_counter[7373] = 4'b0000;
    GSharePlugin_logic_mem_counter[7374] = 4'b0000;
    GSharePlugin_logic_mem_counter[7375] = 4'b0000;
    GSharePlugin_logic_mem_counter[7376] = 4'b0000;
    GSharePlugin_logic_mem_counter[7377] = 4'b0000;
    GSharePlugin_logic_mem_counter[7378] = 4'b0000;
    GSharePlugin_logic_mem_counter[7379] = 4'b0000;
    GSharePlugin_logic_mem_counter[7380] = 4'b0000;
    GSharePlugin_logic_mem_counter[7381] = 4'b0000;
    GSharePlugin_logic_mem_counter[7382] = 4'b0000;
    GSharePlugin_logic_mem_counter[7383] = 4'b0000;
    GSharePlugin_logic_mem_counter[7384] = 4'b0000;
    GSharePlugin_logic_mem_counter[7385] = 4'b0000;
    GSharePlugin_logic_mem_counter[7386] = 4'b0000;
    GSharePlugin_logic_mem_counter[7387] = 4'b0000;
    GSharePlugin_logic_mem_counter[7388] = 4'b0000;
    GSharePlugin_logic_mem_counter[7389] = 4'b0000;
    GSharePlugin_logic_mem_counter[7390] = 4'b0000;
    GSharePlugin_logic_mem_counter[7391] = 4'b0000;
    GSharePlugin_logic_mem_counter[7392] = 4'b0000;
    GSharePlugin_logic_mem_counter[7393] = 4'b0000;
    GSharePlugin_logic_mem_counter[7394] = 4'b0000;
    GSharePlugin_logic_mem_counter[7395] = 4'b0000;
    GSharePlugin_logic_mem_counter[7396] = 4'b0000;
    GSharePlugin_logic_mem_counter[7397] = 4'b0000;
    GSharePlugin_logic_mem_counter[7398] = 4'b0000;
    GSharePlugin_logic_mem_counter[7399] = 4'b0000;
    GSharePlugin_logic_mem_counter[7400] = 4'b0000;
    GSharePlugin_logic_mem_counter[7401] = 4'b0000;
    GSharePlugin_logic_mem_counter[7402] = 4'b0000;
    GSharePlugin_logic_mem_counter[7403] = 4'b0000;
    GSharePlugin_logic_mem_counter[7404] = 4'b0000;
    GSharePlugin_logic_mem_counter[7405] = 4'b0000;
    GSharePlugin_logic_mem_counter[7406] = 4'b0000;
    GSharePlugin_logic_mem_counter[7407] = 4'b0000;
    GSharePlugin_logic_mem_counter[7408] = 4'b0000;
    GSharePlugin_logic_mem_counter[7409] = 4'b0000;
    GSharePlugin_logic_mem_counter[7410] = 4'b0000;
    GSharePlugin_logic_mem_counter[7411] = 4'b0000;
    GSharePlugin_logic_mem_counter[7412] = 4'b0000;
    GSharePlugin_logic_mem_counter[7413] = 4'b0000;
    GSharePlugin_logic_mem_counter[7414] = 4'b0000;
    GSharePlugin_logic_mem_counter[7415] = 4'b0000;
    GSharePlugin_logic_mem_counter[7416] = 4'b0000;
    GSharePlugin_logic_mem_counter[7417] = 4'b0000;
    GSharePlugin_logic_mem_counter[7418] = 4'b0000;
    GSharePlugin_logic_mem_counter[7419] = 4'b0000;
    GSharePlugin_logic_mem_counter[7420] = 4'b0000;
    GSharePlugin_logic_mem_counter[7421] = 4'b0000;
    GSharePlugin_logic_mem_counter[7422] = 4'b0000;
    GSharePlugin_logic_mem_counter[7423] = 4'b0000;
    GSharePlugin_logic_mem_counter[7424] = 4'b0000;
    GSharePlugin_logic_mem_counter[7425] = 4'b0000;
    GSharePlugin_logic_mem_counter[7426] = 4'b0000;
    GSharePlugin_logic_mem_counter[7427] = 4'b0000;
    GSharePlugin_logic_mem_counter[7428] = 4'b0000;
    GSharePlugin_logic_mem_counter[7429] = 4'b0000;
    GSharePlugin_logic_mem_counter[7430] = 4'b0000;
    GSharePlugin_logic_mem_counter[7431] = 4'b0000;
    GSharePlugin_logic_mem_counter[7432] = 4'b0000;
    GSharePlugin_logic_mem_counter[7433] = 4'b0000;
    GSharePlugin_logic_mem_counter[7434] = 4'b0000;
    GSharePlugin_logic_mem_counter[7435] = 4'b0000;
    GSharePlugin_logic_mem_counter[7436] = 4'b0000;
    GSharePlugin_logic_mem_counter[7437] = 4'b0000;
    GSharePlugin_logic_mem_counter[7438] = 4'b0000;
    GSharePlugin_logic_mem_counter[7439] = 4'b0000;
    GSharePlugin_logic_mem_counter[7440] = 4'b0000;
    GSharePlugin_logic_mem_counter[7441] = 4'b0000;
    GSharePlugin_logic_mem_counter[7442] = 4'b0000;
    GSharePlugin_logic_mem_counter[7443] = 4'b0000;
    GSharePlugin_logic_mem_counter[7444] = 4'b0000;
    GSharePlugin_logic_mem_counter[7445] = 4'b0000;
    GSharePlugin_logic_mem_counter[7446] = 4'b0000;
    GSharePlugin_logic_mem_counter[7447] = 4'b0000;
    GSharePlugin_logic_mem_counter[7448] = 4'b0000;
    GSharePlugin_logic_mem_counter[7449] = 4'b0000;
    GSharePlugin_logic_mem_counter[7450] = 4'b0000;
    GSharePlugin_logic_mem_counter[7451] = 4'b0000;
    GSharePlugin_logic_mem_counter[7452] = 4'b0000;
    GSharePlugin_logic_mem_counter[7453] = 4'b0000;
    GSharePlugin_logic_mem_counter[7454] = 4'b0000;
    GSharePlugin_logic_mem_counter[7455] = 4'b0000;
    GSharePlugin_logic_mem_counter[7456] = 4'b0000;
    GSharePlugin_logic_mem_counter[7457] = 4'b0000;
    GSharePlugin_logic_mem_counter[7458] = 4'b0000;
    GSharePlugin_logic_mem_counter[7459] = 4'b0000;
    GSharePlugin_logic_mem_counter[7460] = 4'b0000;
    GSharePlugin_logic_mem_counter[7461] = 4'b0000;
    GSharePlugin_logic_mem_counter[7462] = 4'b0000;
    GSharePlugin_logic_mem_counter[7463] = 4'b0000;
    GSharePlugin_logic_mem_counter[7464] = 4'b0000;
    GSharePlugin_logic_mem_counter[7465] = 4'b0000;
    GSharePlugin_logic_mem_counter[7466] = 4'b0000;
    GSharePlugin_logic_mem_counter[7467] = 4'b0000;
    GSharePlugin_logic_mem_counter[7468] = 4'b0000;
    GSharePlugin_logic_mem_counter[7469] = 4'b0000;
    GSharePlugin_logic_mem_counter[7470] = 4'b0000;
    GSharePlugin_logic_mem_counter[7471] = 4'b0000;
    GSharePlugin_logic_mem_counter[7472] = 4'b0000;
    GSharePlugin_logic_mem_counter[7473] = 4'b0000;
    GSharePlugin_logic_mem_counter[7474] = 4'b0000;
    GSharePlugin_logic_mem_counter[7475] = 4'b0000;
    GSharePlugin_logic_mem_counter[7476] = 4'b0000;
    GSharePlugin_logic_mem_counter[7477] = 4'b0000;
    GSharePlugin_logic_mem_counter[7478] = 4'b0000;
    GSharePlugin_logic_mem_counter[7479] = 4'b0000;
    GSharePlugin_logic_mem_counter[7480] = 4'b0000;
    GSharePlugin_logic_mem_counter[7481] = 4'b0000;
    GSharePlugin_logic_mem_counter[7482] = 4'b0000;
    GSharePlugin_logic_mem_counter[7483] = 4'b0000;
    GSharePlugin_logic_mem_counter[7484] = 4'b0000;
    GSharePlugin_logic_mem_counter[7485] = 4'b0000;
    GSharePlugin_logic_mem_counter[7486] = 4'b0000;
    GSharePlugin_logic_mem_counter[7487] = 4'b0000;
    GSharePlugin_logic_mem_counter[7488] = 4'b0000;
    GSharePlugin_logic_mem_counter[7489] = 4'b0000;
    GSharePlugin_logic_mem_counter[7490] = 4'b0000;
    GSharePlugin_logic_mem_counter[7491] = 4'b0000;
    GSharePlugin_logic_mem_counter[7492] = 4'b0000;
    GSharePlugin_logic_mem_counter[7493] = 4'b0000;
    GSharePlugin_logic_mem_counter[7494] = 4'b0000;
    GSharePlugin_logic_mem_counter[7495] = 4'b0000;
    GSharePlugin_logic_mem_counter[7496] = 4'b0000;
    GSharePlugin_logic_mem_counter[7497] = 4'b0000;
    GSharePlugin_logic_mem_counter[7498] = 4'b0000;
    GSharePlugin_logic_mem_counter[7499] = 4'b0000;
    GSharePlugin_logic_mem_counter[7500] = 4'b0000;
    GSharePlugin_logic_mem_counter[7501] = 4'b0000;
    GSharePlugin_logic_mem_counter[7502] = 4'b0000;
    GSharePlugin_logic_mem_counter[7503] = 4'b0000;
    GSharePlugin_logic_mem_counter[7504] = 4'b0000;
    GSharePlugin_logic_mem_counter[7505] = 4'b0000;
    GSharePlugin_logic_mem_counter[7506] = 4'b0000;
    GSharePlugin_logic_mem_counter[7507] = 4'b0000;
    GSharePlugin_logic_mem_counter[7508] = 4'b0000;
    GSharePlugin_logic_mem_counter[7509] = 4'b0000;
    GSharePlugin_logic_mem_counter[7510] = 4'b0000;
    GSharePlugin_logic_mem_counter[7511] = 4'b0000;
    GSharePlugin_logic_mem_counter[7512] = 4'b0000;
    GSharePlugin_logic_mem_counter[7513] = 4'b0000;
    GSharePlugin_logic_mem_counter[7514] = 4'b0000;
    GSharePlugin_logic_mem_counter[7515] = 4'b0000;
    GSharePlugin_logic_mem_counter[7516] = 4'b0000;
    GSharePlugin_logic_mem_counter[7517] = 4'b0000;
    GSharePlugin_logic_mem_counter[7518] = 4'b0000;
    GSharePlugin_logic_mem_counter[7519] = 4'b0000;
    GSharePlugin_logic_mem_counter[7520] = 4'b0000;
    GSharePlugin_logic_mem_counter[7521] = 4'b0000;
    GSharePlugin_logic_mem_counter[7522] = 4'b0000;
    GSharePlugin_logic_mem_counter[7523] = 4'b0000;
    GSharePlugin_logic_mem_counter[7524] = 4'b0000;
    GSharePlugin_logic_mem_counter[7525] = 4'b0000;
    GSharePlugin_logic_mem_counter[7526] = 4'b0000;
    GSharePlugin_logic_mem_counter[7527] = 4'b0000;
    GSharePlugin_logic_mem_counter[7528] = 4'b0000;
    GSharePlugin_logic_mem_counter[7529] = 4'b0000;
    GSharePlugin_logic_mem_counter[7530] = 4'b0000;
    GSharePlugin_logic_mem_counter[7531] = 4'b0000;
    GSharePlugin_logic_mem_counter[7532] = 4'b0000;
    GSharePlugin_logic_mem_counter[7533] = 4'b0000;
    GSharePlugin_logic_mem_counter[7534] = 4'b0000;
    GSharePlugin_logic_mem_counter[7535] = 4'b0000;
    GSharePlugin_logic_mem_counter[7536] = 4'b0000;
    GSharePlugin_logic_mem_counter[7537] = 4'b0000;
    GSharePlugin_logic_mem_counter[7538] = 4'b0000;
    GSharePlugin_logic_mem_counter[7539] = 4'b0000;
    GSharePlugin_logic_mem_counter[7540] = 4'b0000;
    GSharePlugin_logic_mem_counter[7541] = 4'b0000;
    GSharePlugin_logic_mem_counter[7542] = 4'b0000;
    GSharePlugin_logic_mem_counter[7543] = 4'b0000;
    GSharePlugin_logic_mem_counter[7544] = 4'b0000;
    GSharePlugin_logic_mem_counter[7545] = 4'b0000;
    GSharePlugin_logic_mem_counter[7546] = 4'b0000;
    GSharePlugin_logic_mem_counter[7547] = 4'b0000;
    GSharePlugin_logic_mem_counter[7548] = 4'b0000;
    GSharePlugin_logic_mem_counter[7549] = 4'b0000;
    GSharePlugin_logic_mem_counter[7550] = 4'b0000;
    GSharePlugin_logic_mem_counter[7551] = 4'b0000;
    GSharePlugin_logic_mem_counter[7552] = 4'b0000;
    GSharePlugin_logic_mem_counter[7553] = 4'b0000;
    GSharePlugin_logic_mem_counter[7554] = 4'b0000;
    GSharePlugin_logic_mem_counter[7555] = 4'b0000;
    GSharePlugin_logic_mem_counter[7556] = 4'b0000;
    GSharePlugin_logic_mem_counter[7557] = 4'b0000;
    GSharePlugin_logic_mem_counter[7558] = 4'b0000;
    GSharePlugin_logic_mem_counter[7559] = 4'b0000;
    GSharePlugin_logic_mem_counter[7560] = 4'b0000;
    GSharePlugin_logic_mem_counter[7561] = 4'b0000;
    GSharePlugin_logic_mem_counter[7562] = 4'b0000;
    GSharePlugin_logic_mem_counter[7563] = 4'b0000;
    GSharePlugin_logic_mem_counter[7564] = 4'b0000;
    GSharePlugin_logic_mem_counter[7565] = 4'b0000;
    GSharePlugin_logic_mem_counter[7566] = 4'b0000;
    GSharePlugin_logic_mem_counter[7567] = 4'b0000;
    GSharePlugin_logic_mem_counter[7568] = 4'b0000;
    GSharePlugin_logic_mem_counter[7569] = 4'b0000;
    GSharePlugin_logic_mem_counter[7570] = 4'b0000;
    GSharePlugin_logic_mem_counter[7571] = 4'b0000;
    GSharePlugin_logic_mem_counter[7572] = 4'b0000;
    GSharePlugin_logic_mem_counter[7573] = 4'b0000;
    GSharePlugin_logic_mem_counter[7574] = 4'b0000;
    GSharePlugin_logic_mem_counter[7575] = 4'b0000;
    GSharePlugin_logic_mem_counter[7576] = 4'b0000;
    GSharePlugin_logic_mem_counter[7577] = 4'b0000;
    GSharePlugin_logic_mem_counter[7578] = 4'b0000;
    GSharePlugin_logic_mem_counter[7579] = 4'b0000;
    GSharePlugin_logic_mem_counter[7580] = 4'b0000;
    GSharePlugin_logic_mem_counter[7581] = 4'b0000;
    GSharePlugin_logic_mem_counter[7582] = 4'b0000;
    GSharePlugin_logic_mem_counter[7583] = 4'b0000;
    GSharePlugin_logic_mem_counter[7584] = 4'b0000;
    GSharePlugin_logic_mem_counter[7585] = 4'b0000;
    GSharePlugin_logic_mem_counter[7586] = 4'b0000;
    GSharePlugin_logic_mem_counter[7587] = 4'b0000;
    GSharePlugin_logic_mem_counter[7588] = 4'b0000;
    GSharePlugin_logic_mem_counter[7589] = 4'b0000;
    GSharePlugin_logic_mem_counter[7590] = 4'b0000;
    GSharePlugin_logic_mem_counter[7591] = 4'b0000;
    GSharePlugin_logic_mem_counter[7592] = 4'b0000;
    GSharePlugin_logic_mem_counter[7593] = 4'b0000;
    GSharePlugin_logic_mem_counter[7594] = 4'b0000;
    GSharePlugin_logic_mem_counter[7595] = 4'b0000;
    GSharePlugin_logic_mem_counter[7596] = 4'b0000;
    GSharePlugin_logic_mem_counter[7597] = 4'b0000;
    GSharePlugin_logic_mem_counter[7598] = 4'b0000;
    GSharePlugin_logic_mem_counter[7599] = 4'b0000;
    GSharePlugin_logic_mem_counter[7600] = 4'b0000;
    GSharePlugin_logic_mem_counter[7601] = 4'b0000;
    GSharePlugin_logic_mem_counter[7602] = 4'b0000;
    GSharePlugin_logic_mem_counter[7603] = 4'b0000;
    GSharePlugin_logic_mem_counter[7604] = 4'b0000;
    GSharePlugin_logic_mem_counter[7605] = 4'b0000;
    GSharePlugin_logic_mem_counter[7606] = 4'b0000;
    GSharePlugin_logic_mem_counter[7607] = 4'b0000;
    GSharePlugin_logic_mem_counter[7608] = 4'b0000;
    GSharePlugin_logic_mem_counter[7609] = 4'b0000;
    GSharePlugin_logic_mem_counter[7610] = 4'b0000;
    GSharePlugin_logic_mem_counter[7611] = 4'b0000;
    GSharePlugin_logic_mem_counter[7612] = 4'b0000;
    GSharePlugin_logic_mem_counter[7613] = 4'b0000;
    GSharePlugin_logic_mem_counter[7614] = 4'b0000;
    GSharePlugin_logic_mem_counter[7615] = 4'b0000;
    GSharePlugin_logic_mem_counter[7616] = 4'b0000;
    GSharePlugin_logic_mem_counter[7617] = 4'b0000;
    GSharePlugin_logic_mem_counter[7618] = 4'b0000;
    GSharePlugin_logic_mem_counter[7619] = 4'b0000;
    GSharePlugin_logic_mem_counter[7620] = 4'b0000;
    GSharePlugin_logic_mem_counter[7621] = 4'b0000;
    GSharePlugin_logic_mem_counter[7622] = 4'b0000;
    GSharePlugin_logic_mem_counter[7623] = 4'b0000;
    GSharePlugin_logic_mem_counter[7624] = 4'b0000;
    GSharePlugin_logic_mem_counter[7625] = 4'b0000;
    GSharePlugin_logic_mem_counter[7626] = 4'b0000;
    GSharePlugin_logic_mem_counter[7627] = 4'b0000;
    GSharePlugin_logic_mem_counter[7628] = 4'b0000;
    GSharePlugin_logic_mem_counter[7629] = 4'b0000;
    GSharePlugin_logic_mem_counter[7630] = 4'b0000;
    GSharePlugin_logic_mem_counter[7631] = 4'b0000;
    GSharePlugin_logic_mem_counter[7632] = 4'b0000;
    GSharePlugin_logic_mem_counter[7633] = 4'b0000;
    GSharePlugin_logic_mem_counter[7634] = 4'b0000;
    GSharePlugin_logic_mem_counter[7635] = 4'b0000;
    GSharePlugin_logic_mem_counter[7636] = 4'b0000;
    GSharePlugin_logic_mem_counter[7637] = 4'b0000;
    GSharePlugin_logic_mem_counter[7638] = 4'b0000;
    GSharePlugin_logic_mem_counter[7639] = 4'b0000;
    GSharePlugin_logic_mem_counter[7640] = 4'b0000;
    GSharePlugin_logic_mem_counter[7641] = 4'b0000;
    GSharePlugin_logic_mem_counter[7642] = 4'b0000;
    GSharePlugin_logic_mem_counter[7643] = 4'b0000;
    GSharePlugin_logic_mem_counter[7644] = 4'b0000;
    GSharePlugin_logic_mem_counter[7645] = 4'b0000;
    GSharePlugin_logic_mem_counter[7646] = 4'b0000;
    GSharePlugin_logic_mem_counter[7647] = 4'b0000;
    GSharePlugin_logic_mem_counter[7648] = 4'b0000;
    GSharePlugin_logic_mem_counter[7649] = 4'b0000;
    GSharePlugin_logic_mem_counter[7650] = 4'b0000;
    GSharePlugin_logic_mem_counter[7651] = 4'b0000;
    GSharePlugin_logic_mem_counter[7652] = 4'b0000;
    GSharePlugin_logic_mem_counter[7653] = 4'b0000;
    GSharePlugin_logic_mem_counter[7654] = 4'b0000;
    GSharePlugin_logic_mem_counter[7655] = 4'b0000;
    GSharePlugin_logic_mem_counter[7656] = 4'b0000;
    GSharePlugin_logic_mem_counter[7657] = 4'b0000;
    GSharePlugin_logic_mem_counter[7658] = 4'b0000;
    GSharePlugin_logic_mem_counter[7659] = 4'b0000;
    GSharePlugin_logic_mem_counter[7660] = 4'b0000;
    GSharePlugin_logic_mem_counter[7661] = 4'b0000;
    GSharePlugin_logic_mem_counter[7662] = 4'b0000;
    GSharePlugin_logic_mem_counter[7663] = 4'b0000;
    GSharePlugin_logic_mem_counter[7664] = 4'b0000;
    GSharePlugin_logic_mem_counter[7665] = 4'b0000;
    GSharePlugin_logic_mem_counter[7666] = 4'b0000;
    GSharePlugin_logic_mem_counter[7667] = 4'b0000;
    GSharePlugin_logic_mem_counter[7668] = 4'b0000;
    GSharePlugin_logic_mem_counter[7669] = 4'b0000;
    GSharePlugin_logic_mem_counter[7670] = 4'b0000;
    GSharePlugin_logic_mem_counter[7671] = 4'b0000;
    GSharePlugin_logic_mem_counter[7672] = 4'b0000;
    GSharePlugin_logic_mem_counter[7673] = 4'b0000;
    GSharePlugin_logic_mem_counter[7674] = 4'b0000;
    GSharePlugin_logic_mem_counter[7675] = 4'b0000;
    GSharePlugin_logic_mem_counter[7676] = 4'b0000;
    GSharePlugin_logic_mem_counter[7677] = 4'b0000;
    GSharePlugin_logic_mem_counter[7678] = 4'b0000;
    GSharePlugin_logic_mem_counter[7679] = 4'b0000;
    GSharePlugin_logic_mem_counter[7680] = 4'b0000;
    GSharePlugin_logic_mem_counter[7681] = 4'b0000;
    GSharePlugin_logic_mem_counter[7682] = 4'b0000;
    GSharePlugin_logic_mem_counter[7683] = 4'b0000;
    GSharePlugin_logic_mem_counter[7684] = 4'b0000;
    GSharePlugin_logic_mem_counter[7685] = 4'b0000;
    GSharePlugin_logic_mem_counter[7686] = 4'b0000;
    GSharePlugin_logic_mem_counter[7687] = 4'b0000;
    GSharePlugin_logic_mem_counter[7688] = 4'b0000;
    GSharePlugin_logic_mem_counter[7689] = 4'b0000;
    GSharePlugin_logic_mem_counter[7690] = 4'b0000;
    GSharePlugin_logic_mem_counter[7691] = 4'b0000;
    GSharePlugin_logic_mem_counter[7692] = 4'b0000;
    GSharePlugin_logic_mem_counter[7693] = 4'b0000;
    GSharePlugin_logic_mem_counter[7694] = 4'b0000;
    GSharePlugin_logic_mem_counter[7695] = 4'b0000;
    GSharePlugin_logic_mem_counter[7696] = 4'b0000;
    GSharePlugin_logic_mem_counter[7697] = 4'b0000;
    GSharePlugin_logic_mem_counter[7698] = 4'b0000;
    GSharePlugin_logic_mem_counter[7699] = 4'b0000;
    GSharePlugin_logic_mem_counter[7700] = 4'b0000;
    GSharePlugin_logic_mem_counter[7701] = 4'b0000;
    GSharePlugin_logic_mem_counter[7702] = 4'b0000;
    GSharePlugin_logic_mem_counter[7703] = 4'b0000;
    GSharePlugin_logic_mem_counter[7704] = 4'b0000;
    GSharePlugin_logic_mem_counter[7705] = 4'b0000;
    GSharePlugin_logic_mem_counter[7706] = 4'b0000;
    GSharePlugin_logic_mem_counter[7707] = 4'b0000;
    GSharePlugin_logic_mem_counter[7708] = 4'b0000;
    GSharePlugin_logic_mem_counter[7709] = 4'b0000;
    GSharePlugin_logic_mem_counter[7710] = 4'b0000;
    GSharePlugin_logic_mem_counter[7711] = 4'b0000;
    GSharePlugin_logic_mem_counter[7712] = 4'b0000;
    GSharePlugin_logic_mem_counter[7713] = 4'b0000;
    GSharePlugin_logic_mem_counter[7714] = 4'b0000;
    GSharePlugin_logic_mem_counter[7715] = 4'b0000;
    GSharePlugin_logic_mem_counter[7716] = 4'b0000;
    GSharePlugin_logic_mem_counter[7717] = 4'b0000;
    GSharePlugin_logic_mem_counter[7718] = 4'b0000;
    GSharePlugin_logic_mem_counter[7719] = 4'b0000;
    GSharePlugin_logic_mem_counter[7720] = 4'b0000;
    GSharePlugin_logic_mem_counter[7721] = 4'b0000;
    GSharePlugin_logic_mem_counter[7722] = 4'b0000;
    GSharePlugin_logic_mem_counter[7723] = 4'b0000;
    GSharePlugin_logic_mem_counter[7724] = 4'b0000;
    GSharePlugin_logic_mem_counter[7725] = 4'b0000;
    GSharePlugin_logic_mem_counter[7726] = 4'b0000;
    GSharePlugin_logic_mem_counter[7727] = 4'b0000;
    GSharePlugin_logic_mem_counter[7728] = 4'b0000;
    GSharePlugin_logic_mem_counter[7729] = 4'b0000;
    GSharePlugin_logic_mem_counter[7730] = 4'b0000;
    GSharePlugin_logic_mem_counter[7731] = 4'b0000;
    GSharePlugin_logic_mem_counter[7732] = 4'b0000;
    GSharePlugin_logic_mem_counter[7733] = 4'b0000;
    GSharePlugin_logic_mem_counter[7734] = 4'b0000;
    GSharePlugin_logic_mem_counter[7735] = 4'b0000;
    GSharePlugin_logic_mem_counter[7736] = 4'b0000;
    GSharePlugin_logic_mem_counter[7737] = 4'b0000;
    GSharePlugin_logic_mem_counter[7738] = 4'b0000;
    GSharePlugin_logic_mem_counter[7739] = 4'b0000;
    GSharePlugin_logic_mem_counter[7740] = 4'b0000;
    GSharePlugin_logic_mem_counter[7741] = 4'b0000;
    GSharePlugin_logic_mem_counter[7742] = 4'b0000;
    GSharePlugin_logic_mem_counter[7743] = 4'b0000;
    GSharePlugin_logic_mem_counter[7744] = 4'b0000;
    GSharePlugin_logic_mem_counter[7745] = 4'b0000;
    GSharePlugin_logic_mem_counter[7746] = 4'b0000;
    GSharePlugin_logic_mem_counter[7747] = 4'b0000;
    GSharePlugin_logic_mem_counter[7748] = 4'b0000;
    GSharePlugin_logic_mem_counter[7749] = 4'b0000;
    GSharePlugin_logic_mem_counter[7750] = 4'b0000;
    GSharePlugin_logic_mem_counter[7751] = 4'b0000;
    GSharePlugin_logic_mem_counter[7752] = 4'b0000;
    GSharePlugin_logic_mem_counter[7753] = 4'b0000;
    GSharePlugin_logic_mem_counter[7754] = 4'b0000;
    GSharePlugin_logic_mem_counter[7755] = 4'b0000;
    GSharePlugin_logic_mem_counter[7756] = 4'b0000;
    GSharePlugin_logic_mem_counter[7757] = 4'b0000;
    GSharePlugin_logic_mem_counter[7758] = 4'b0000;
    GSharePlugin_logic_mem_counter[7759] = 4'b0000;
    GSharePlugin_logic_mem_counter[7760] = 4'b0000;
    GSharePlugin_logic_mem_counter[7761] = 4'b0000;
    GSharePlugin_logic_mem_counter[7762] = 4'b0000;
    GSharePlugin_logic_mem_counter[7763] = 4'b0000;
    GSharePlugin_logic_mem_counter[7764] = 4'b0000;
    GSharePlugin_logic_mem_counter[7765] = 4'b0000;
    GSharePlugin_logic_mem_counter[7766] = 4'b0000;
    GSharePlugin_logic_mem_counter[7767] = 4'b0000;
    GSharePlugin_logic_mem_counter[7768] = 4'b0000;
    GSharePlugin_logic_mem_counter[7769] = 4'b0000;
    GSharePlugin_logic_mem_counter[7770] = 4'b0000;
    GSharePlugin_logic_mem_counter[7771] = 4'b0000;
    GSharePlugin_logic_mem_counter[7772] = 4'b0000;
    GSharePlugin_logic_mem_counter[7773] = 4'b0000;
    GSharePlugin_logic_mem_counter[7774] = 4'b0000;
    GSharePlugin_logic_mem_counter[7775] = 4'b0000;
    GSharePlugin_logic_mem_counter[7776] = 4'b0000;
    GSharePlugin_logic_mem_counter[7777] = 4'b0000;
    GSharePlugin_logic_mem_counter[7778] = 4'b0000;
    GSharePlugin_logic_mem_counter[7779] = 4'b0000;
    GSharePlugin_logic_mem_counter[7780] = 4'b0000;
    GSharePlugin_logic_mem_counter[7781] = 4'b0000;
    GSharePlugin_logic_mem_counter[7782] = 4'b0000;
    GSharePlugin_logic_mem_counter[7783] = 4'b0000;
    GSharePlugin_logic_mem_counter[7784] = 4'b0000;
    GSharePlugin_logic_mem_counter[7785] = 4'b0000;
    GSharePlugin_logic_mem_counter[7786] = 4'b0000;
    GSharePlugin_logic_mem_counter[7787] = 4'b0000;
    GSharePlugin_logic_mem_counter[7788] = 4'b0000;
    GSharePlugin_logic_mem_counter[7789] = 4'b0000;
    GSharePlugin_logic_mem_counter[7790] = 4'b0000;
    GSharePlugin_logic_mem_counter[7791] = 4'b0000;
    GSharePlugin_logic_mem_counter[7792] = 4'b0000;
    GSharePlugin_logic_mem_counter[7793] = 4'b0000;
    GSharePlugin_logic_mem_counter[7794] = 4'b0000;
    GSharePlugin_logic_mem_counter[7795] = 4'b0000;
    GSharePlugin_logic_mem_counter[7796] = 4'b0000;
    GSharePlugin_logic_mem_counter[7797] = 4'b0000;
    GSharePlugin_logic_mem_counter[7798] = 4'b0000;
    GSharePlugin_logic_mem_counter[7799] = 4'b0000;
    GSharePlugin_logic_mem_counter[7800] = 4'b0000;
    GSharePlugin_logic_mem_counter[7801] = 4'b0000;
    GSharePlugin_logic_mem_counter[7802] = 4'b0000;
    GSharePlugin_logic_mem_counter[7803] = 4'b0000;
    GSharePlugin_logic_mem_counter[7804] = 4'b0000;
    GSharePlugin_logic_mem_counter[7805] = 4'b0000;
    GSharePlugin_logic_mem_counter[7806] = 4'b0000;
    GSharePlugin_logic_mem_counter[7807] = 4'b0000;
    GSharePlugin_logic_mem_counter[7808] = 4'b0000;
    GSharePlugin_logic_mem_counter[7809] = 4'b0000;
    GSharePlugin_logic_mem_counter[7810] = 4'b0000;
    GSharePlugin_logic_mem_counter[7811] = 4'b0000;
    GSharePlugin_logic_mem_counter[7812] = 4'b0000;
    GSharePlugin_logic_mem_counter[7813] = 4'b0000;
    GSharePlugin_logic_mem_counter[7814] = 4'b0000;
    GSharePlugin_logic_mem_counter[7815] = 4'b0000;
    GSharePlugin_logic_mem_counter[7816] = 4'b0000;
    GSharePlugin_logic_mem_counter[7817] = 4'b0000;
    GSharePlugin_logic_mem_counter[7818] = 4'b0000;
    GSharePlugin_logic_mem_counter[7819] = 4'b0000;
    GSharePlugin_logic_mem_counter[7820] = 4'b0000;
    GSharePlugin_logic_mem_counter[7821] = 4'b0000;
    GSharePlugin_logic_mem_counter[7822] = 4'b0000;
    GSharePlugin_logic_mem_counter[7823] = 4'b0000;
    GSharePlugin_logic_mem_counter[7824] = 4'b0000;
    GSharePlugin_logic_mem_counter[7825] = 4'b0000;
    GSharePlugin_logic_mem_counter[7826] = 4'b0000;
    GSharePlugin_logic_mem_counter[7827] = 4'b0000;
    GSharePlugin_logic_mem_counter[7828] = 4'b0000;
    GSharePlugin_logic_mem_counter[7829] = 4'b0000;
    GSharePlugin_logic_mem_counter[7830] = 4'b0000;
    GSharePlugin_logic_mem_counter[7831] = 4'b0000;
    GSharePlugin_logic_mem_counter[7832] = 4'b0000;
    GSharePlugin_logic_mem_counter[7833] = 4'b0000;
    GSharePlugin_logic_mem_counter[7834] = 4'b0000;
    GSharePlugin_logic_mem_counter[7835] = 4'b0000;
    GSharePlugin_logic_mem_counter[7836] = 4'b0000;
    GSharePlugin_logic_mem_counter[7837] = 4'b0000;
    GSharePlugin_logic_mem_counter[7838] = 4'b0000;
    GSharePlugin_logic_mem_counter[7839] = 4'b0000;
    GSharePlugin_logic_mem_counter[7840] = 4'b0000;
    GSharePlugin_logic_mem_counter[7841] = 4'b0000;
    GSharePlugin_logic_mem_counter[7842] = 4'b0000;
    GSharePlugin_logic_mem_counter[7843] = 4'b0000;
    GSharePlugin_logic_mem_counter[7844] = 4'b0000;
    GSharePlugin_logic_mem_counter[7845] = 4'b0000;
    GSharePlugin_logic_mem_counter[7846] = 4'b0000;
    GSharePlugin_logic_mem_counter[7847] = 4'b0000;
    GSharePlugin_logic_mem_counter[7848] = 4'b0000;
    GSharePlugin_logic_mem_counter[7849] = 4'b0000;
    GSharePlugin_logic_mem_counter[7850] = 4'b0000;
    GSharePlugin_logic_mem_counter[7851] = 4'b0000;
    GSharePlugin_logic_mem_counter[7852] = 4'b0000;
    GSharePlugin_logic_mem_counter[7853] = 4'b0000;
    GSharePlugin_logic_mem_counter[7854] = 4'b0000;
    GSharePlugin_logic_mem_counter[7855] = 4'b0000;
    GSharePlugin_logic_mem_counter[7856] = 4'b0000;
    GSharePlugin_logic_mem_counter[7857] = 4'b0000;
    GSharePlugin_logic_mem_counter[7858] = 4'b0000;
    GSharePlugin_logic_mem_counter[7859] = 4'b0000;
    GSharePlugin_logic_mem_counter[7860] = 4'b0000;
    GSharePlugin_logic_mem_counter[7861] = 4'b0000;
    GSharePlugin_logic_mem_counter[7862] = 4'b0000;
    GSharePlugin_logic_mem_counter[7863] = 4'b0000;
    GSharePlugin_logic_mem_counter[7864] = 4'b0000;
    GSharePlugin_logic_mem_counter[7865] = 4'b0000;
    GSharePlugin_logic_mem_counter[7866] = 4'b0000;
    GSharePlugin_logic_mem_counter[7867] = 4'b0000;
    GSharePlugin_logic_mem_counter[7868] = 4'b0000;
    GSharePlugin_logic_mem_counter[7869] = 4'b0000;
    GSharePlugin_logic_mem_counter[7870] = 4'b0000;
    GSharePlugin_logic_mem_counter[7871] = 4'b0000;
    GSharePlugin_logic_mem_counter[7872] = 4'b0000;
    GSharePlugin_logic_mem_counter[7873] = 4'b0000;
    GSharePlugin_logic_mem_counter[7874] = 4'b0000;
    GSharePlugin_logic_mem_counter[7875] = 4'b0000;
    GSharePlugin_logic_mem_counter[7876] = 4'b0000;
    GSharePlugin_logic_mem_counter[7877] = 4'b0000;
    GSharePlugin_logic_mem_counter[7878] = 4'b0000;
    GSharePlugin_logic_mem_counter[7879] = 4'b0000;
    GSharePlugin_logic_mem_counter[7880] = 4'b0000;
    GSharePlugin_logic_mem_counter[7881] = 4'b0000;
    GSharePlugin_logic_mem_counter[7882] = 4'b0000;
    GSharePlugin_logic_mem_counter[7883] = 4'b0000;
    GSharePlugin_logic_mem_counter[7884] = 4'b0000;
    GSharePlugin_logic_mem_counter[7885] = 4'b0000;
    GSharePlugin_logic_mem_counter[7886] = 4'b0000;
    GSharePlugin_logic_mem_counter[7887] = 4'b0000;
    GSharePlugin_logic_mem_counter[7888] = 4'b0000;
    GSharePlugin_logic_mem_counter[7889] = 4'b0000;
    GSharePlugin_logic_mem_counter[7890] = 4'b0000;
    GSharePlugin_logic_mem_counter[7891] = 4'b0000;
    GSharePlugin_logic_mem_counter[7892] = 4'b0000;
    GSharePlugin_logic_mem_counter[7893] = 4'b0000;
    GSharePlugin_logic_mem_counter[7894] = 4'b0000;
    GSharePlugin_logic_mem_counter[7895] = 4'b0000;
    GSharePlugin_logic_mem_counter[7896] = 4'b0000;
    GSharePlugin_logic_mem_counter[7897] = 4'b0000;
    GSharePlugin_logic_mem_counter[7898] = 4'b0000;
    GSharePlugin_logic_mem_counter[7899] = 4'b0000;
    GSharePlugin_logic_mem_counter[7900] = 4'b0000;
    GSharePlugin_logic_mem_counter[7901] = 4'b0000;
    GSharePlugin_logic_mem_counter[7902] = 4'b0000;
    GSharePlugin_logic_mem_counter[7903] = 4'b0000;
    GSharePlugin_logic_mem_counter[7904] = 4'b0000;
    GSharePlugin_logic_mem_counter[7905] = 4'b0000;
    GSharePlugin_logic_mem_counter[7906] = 4'b0000;
    GSharePlugin_logic_mem_counter[7907] = 4'b0000;
    GSharePlugin_logic_mem_counter[7908] = 4'b0000;
    GSharePlugin_logic_mem_counter[7909] = 4'b0000;
    GSharePlugin_logic_mem_counter[7910] = 4'b0000;
    GSharePlugin_logic_mem_counter[7911] = 4'b0000;
    GSharePlugin_logic_mem_counter[7912] = 4'b0000;
    GSharePlugin_logic_mem_counter[7913] = 4'b0000;
    GSharePlugin_logic_mem_counter[7914] = 4'b0000;
    GSharePlugin_logic_mem_counter[7915] = 4'b0000;
    GSharePlugin_logic_mem_counter[7916] = 4'b0000;
    GSharePlugin_logic_mem_counter[7917] = 4'b0000;
    GSharePlugin_logic_mem_counter[7918] = 4'b0000;
    GSharePlugin_logic_mem_counter[7919] = 4'b0000;
    GSharePlugin_logic_mem_counter[7920] = 4'b0000;
    GSharePlugin_logic_mem_counter[7921] = 4'b0000;
    GSharePlugin_logic_mem_counter[7922] = 4'b0000;
    GSharePlugin_logic_mem_counter[7923] = 4'b0000;
    GSharePlugin_logic_mem_counter[7924] = 4'b0000;
    GSharePlugin_logic_mem_counter[7925] = 4'b0000;
    GSharePlugin_logic_mem_counter[7926] = 4'b0000;
    GSharePlugin_logic_mem_counter[7927] = 4'b0000;
    GSharePlugin_logic_mem_counter[7928] = 4'b0000;
    GSharePlugin_logic_mem_counter[7929] = 4'b0000;
    GSharePlugin_logic_mem_counter[7930] = 4'b0000;
    GSharePlugin_logic_mem_counter[7931] = 4'b0000;
    GSharePlugin_logic_mem_counter[7932] = 4'b0000;
    GSharePlugin_logic_mem_counter[7933] = 4'b0000;
    GSharePlugin_logic_mem_counter[7934] = 4'b0000;
    GSharePlugin_logic_mem_counter[7935] = 4'b0000;
    GSharePlugin_logic_mem_counter[7936] = 4'b0000;
    GSharePlugin_logic_mem_counter[7937] = 4'b0000;
    GSharePlugin_logic_mem_counter[7938] = 4'b0000;
    GSharePlugin_logic_mem_counter[7939] = 4'b0000;
    GSharePlugin_logic_mem_counter[7940] = 4'b0000;
    GSharePlugin_logic_mem_counter[7941] = 4'b0000;
    GSharePlugin_logic_mem_counter[7942] = 4'b0000;
    GSharePlugin_logic_mem_counter[7943] = 4'b0000;
    GSharePlugin_logic_mem_counter[7944] = 4'b0000;
    GSharePlugin_logic_mem_counter[7945] = 4'b0000;
    GSharePlugin_logic_mem_counter[7946] = 4'b0000;
    GSharePlugin_logic_mem_counter[7947] = 4'b0000;
    GSharePlugin_logic_mem_counter[7948] = 4'b0000;
    GSharePlugin_logic_mem_counter[7949] = 4'b0000;
    GSharePlugin_logic_mem_counter[7950] = 4'b0000;
    GSharePlugin_logic_mem_counter[7951] = 4'b0000;
    GSharePlugin_logic_mem_counter[7952] = 4'b0000;
    GSharePlugin_logic_mem_counter[7953] = 4'b0000;
    GSharePlugin_logic_mem_counter[7954] = 4'b0000;
    GSharePlugin_logic_mem_counter[7955] = 4'b0000;
    GSharePlugin_logic_mem_counter[7956] = 4'b0000;
    GSharePlugin_logic_mem_counter[7957] = 4'b0000;
    GSharePlugin_logic_mem_counter[7958] = 4'b0000;
    GSharePlugin_logic_mem_counter[7959] = 4'b0000;
    GSharePlugin_logic_mem_counter[7960] = 4'b0000;
    GSharePlugin_logic_mem_counter[7961] = 4'b0000;
    GSharePlugin_logic_mem_counter[7962] = 4'b0000;
    GSharePlugin_logic_mem_counter[7963] = 4'b0000;
    GSharePlugin_logic_mem_counter[7964] = 4'b0000;
    GSharePlugin_logic_mem_counter[7965] = 4'b0000;
    GSharePlugin_logic_mem_counter[7966] = 4'b0000;
    GSharePlugin_logic_mem_counter[7967] = 4'b0000;
    GSharePlugin_logic_mem_counter[7968] = 4'b0000;
    GSharePlugin_logic_mem_counter[7969] = 4'b0000;
    GSharePlugin_logic_mem_counter[7970] = 4'b0000;
    GSharePlugin_logic_mem_counter[7971] = 4'b0000;
    GSharePlugin_logic_mem_counter[7972] = 4'b0000;
    GSharePlugin_logic_mem_counter[7973] = 4'b0000;
    GSharePlugin_logic_mem_counter[7974] = 4'b0000;
    GSharePlugin_logic_mem_counter[7975] = 4'b0000;
    GSharePlugin_logic_mem_counter[7976] = 4'b0000;
    GSharePlugin_logic_mem_counter[7977] = 4'b0000;
    GSharePlugin_logic_mem_counter[7978] = 4'b0000;
    GSharePlugin_logic_mem_counter[7979] = 4'b0000;
    GSharePlugin_logic_mem_counter[7980] = 4'b0000;
    GSharePlugin_logic_mem_counter[7981] = 4'b0000;
    GSharePlugin_logic_mem_counter[7982] = 4'b0000;
    GSharePlugin_logic_mem_counter[7983] = 4'b0000;
    GSharePlugin_logic_mem_counter[7984] = 4'b0000;
    GSharePlugin_logic_mem_counter[7985] = 4'b0000;
    GSharePlugin_logic_mem_counter[7986] = 4'b0000;
    GSharePlugin_logic_mem_counter[7987] = 4'b0000;
    GSharePlugin_logic_mem_counter[7988] = 4'b0000;
    GSharePlugin_logic_mem_counter[7989] = 4'b0000;
    GSharePlugin_logic_mem_counter[7990] = 4'b0000;
    GSharePlugin_logic_mem_counter[7991] = 4'b0000;
    GSharePlugin_logic_mem_counter[7992] = 4'b0000;
    GSharePlugin_logic_mem_counter[7993] = 4'b0000;
    GSharePlugin_logic_mem_counter[7994] = 4'b0000;
    GSharePlugin_logic_mem_counter[7995] = 4'b0000;
    GSharePlugin_logic_mem_counter[7996] = 4'b0000;
    GSharePlugin_logic_mem_counter[7997] = 4'b0000;
    GSharePlugin_logic_mem_counter[7998] = 4'b0000;
    GSharePlugin_logic_mem_counter[7999] = 4'b0000;
    GSharePlugin_logic_mem_counter[8000] = 4'b0000;
    GSharePlugin_logic_mem_counter[8001] = 4'b0000;
    GSharePlugin_logic_mem_counter[8002] = 4'b0000;
    GSharePlugin_logic_mem_counter[8003] = 4'b0000;
    GSharePlugin_logic_mem_counter[8004] = 4'b0000;
    GSharePlugin_logic_mem_counter[8005] = 4'b0000;
    GSharePlugin_logic_mem_counter[8006] = 4'b0000;
    GSharePlugin_logic_mem_counter[8007] = 4'b0000;
    GSharePlugin_logic_mem_counter[8008] = 4'b0000;
    GSharePlugin_logic_mem_counter[8009] = 4'b0000;
    GSharePlugin_logic_mem_counter[8010] = 4'b0000;
    GSharePlugin_logic_mem_counter[8011] = 4'b0000;
    GSharePlugin_logic_mem_counter[8012] = 4'b0000;
    GSharePlugin_logic_mem_counter[8013] = 4'b0000;
    GSharePlugin_logic_mem_counter[8014] = 4'b0000;
    GSharePlugin_logic_mem_counter[8015] = 4'b0000;
    GSharePlugin_logic_mem_counter[8016] = 4'b0000;
    GSharePlugin_logic_mem_counter[8017] = 4'b0000;
    GSharePlugin_logic_mem_counter[8018] = 4'b0000;
    GSharePlugin_logic_mem_counter[8019] = 4'b0000;
    GSharePlugin_logic_mem_counter[8020] = 4'b0000;
    GSharePlugin_logic_mem_counter[8021] = 4'b0000;
    GSharePlugin_logic_mem_counter[8022] = 4'b0000;
    GSharePlugin_logic_mem_counter[8023] = 4'b0000;
    GSharePlugin_logic_mem_counter[8024] = 4'b0000;
    GSharePlugin_logic_mem_counter[8025] = 4'b0000;
    GSharePlugin_logic_mem_counter[8026] = 4'b0000;
    GSharePlugin_logic_mem_counter[8027] = 4'b0000;
    GSharePlugin_logic_mem_counter[8028] = 4'b0000;
    GSharePlugin_logic_mem_counter[8029] = 4'b0000;
    GSharePlugin_logic_mem_counter[8030] = 4'b0000;
    GSharePlugin_logic_mem_counter[8031] = 4'b0000;
    GSharePlugin_logic_mem_counter[8032] = 4'b0000;
    GSharePlugin_logic_mem_counter[8033] = 4'b0000;
    GSharePlugin_logic_mem_counter[8034] = 4'b0000;
    GSharePlugin_logic_mem_counter[8035] = 4'b0000;
    GSharePlugin_logic_mem_counter[8036] = 4'b0000;
    GSharePlugin_logic_mem_counter[8037] = 4'b0000;
    GSharePlugin_logic_mem_counter[8038] = 4'b0000;
    GSharePlugin_logic_mem_counter[8039] = 4'b0000;
    GSharePlugin_logic_mem_counter[8040] = 4'b0000;
    GSharePlugin_logic_mem_counter[8041] = 4'b0000;
    GSharePlugin_logic_mem_counter[8042] = 4'b0000;
    GSharePlugin_logic_mem_counter[8043] = 4'b0000;
    GSharePlugin_logic_mem_counter[8044] = 4'b0000;
    GSharePlugin_logic_mem_counter[8045] = 4'b0000;
    GSharePlugin_logic_mem_counter[8046] = 4'b0000;
    GSharePlugin_logic_mem_counter[8047] = 4'b0000;
    GSharePlugin_logic_mem_counter[8048] = 4'b0000;
    GSharePlugin_logic_mem_counter[8049] = 4'b0000;
    GSharePlugin_logic_mem_counter[8050] = 4'b0000;
    GSharePlugin_logic_mem_counter[8051] = 4'b0000;
    GSharePlugin_logic_mem_counter[8052] = 4'b0000;
    GSharePlugin_logic_mem_counter[8053] = 4'b0000;
    GSharePlugin_logic_mem_counter[8054] = 4'b0000;
    GSharePlugin_logic_mem_counter[8055] = 4'b0000;
    GSharePlugin_logic_mem_counter[8056] = 4'b0000;
    GSharePlugin_logic_mem_counter[8057] = 4'b0000;
    GSharePlugin_logic_mem_counter[8058] = 4'b0000;
    GSharePlugin_logic_mem_counter[8059] = 4'b0000;
    GSharePlugin_logic_mem_counter[8060] = 4'b0000;
    GSharePlugin_logic_mem_counter[8061] = 4'b0000;
    GSharePlugin_logic_mem_counter[8062] = 4'b0000;
    GSharePlugin_logic_mem_counter[8063] = 4'b0000;
    GSharePlugin_logic_mem_counter[8064] = 4'b0000;
    GSharePlugin_logic_mem_counter[8065] = 4'b0000;
    GSharePlugin_logic_mem_counter[8066] = 4'b0000;
    GSharePlugin_logic_mem_counter[8067] = 4'b0000;
    GSharePlugin_logic_mem_counter[8068] = 4'b0000;
    GSharePlugin_logic_mem_counter[8069] = 4'b0000;
    GSharePlugin_logic_mem_counter[8070] = 4'b0000;
    GSharePlugin_logic_mem_counter[8071] = 4'b0000;
    GSharePlugin_logic_mem_counter[8072] = 4'b0000;
    GSharePlugin_logic_mem_counter[8073] = 4'b0000;
    GSharePlugin_logic_mem_counter[8074] = 4'b0000;
    GSharePlugin_logic_mem_counter[8075] = 4'b0000;
    GSharePlugin_logic_mem_counter[8076] = 4'b0000;
    GSharePlugin_logic_mem_counter[8077] = 4'b0000;
    GSharePlugin_logic_mem_counter[8078] = 4'b0000;
    GSharePlugin_logic_mem_counter[8079] = 4'b0000;
    GSharePlugin_logic_mem_counter[8080] = 4'b0000;
    GSharePlugin_logic_mem_counter[8081] = 4'b0000;
    GSharePlugin_logic_mem_counter[8082] = 4'b0000;
    GSharePlugin_logic_mem_counter[8083] = 4'b0000;
    GSharePlugin_logic_mem_counter[8084] = 4'b0000;
    GSharePlugin_logic_mem_counter[8085] = 4'b0000;
    GSharePlugin_logic_mem_counter[8086] = 4'b0000;
    GSharePlugin_logic_mem_counter[8087] = 4'b0000;
    GSharePlugin_logic_mem_counter[8088] = 4'b0000;
    GSharePlugin_logic_mem_counter[8089] = 4'b0000;
    GSharePlugin_logic_mem_counter[8090] = 4'b0000;
    GSharePlugin_logic_mem_counter[8091] = 4'b0000;
    GSharePlugin_logic_mem_counter[8092] = 4'b0000;
    GSharePlugin_logic_mem_counter[8093] = 4'b0000;
    GSharePlugin_logic_mem_counter[8094] = 4'b0000;
    GSharePlugin_logic_mem_counter[8095] = 4'b0000;
    GSharePlugin_logic_mem_counter[8096] = 4'b0000;
    GSharePlugin_logic_mem_counter[8097] = 4'b0000;
    GSharePlugin_logic_mem_counter[8098] = 4'b0000;
    GSharePlugin_logic_mem_counter[8099] = 4'b0000;
    GSharePlugin_logic_mem_counter[8100] = 4'b0000;
    GSharePlugin_logic_mem_counter[8101] = 4'b0000;
    GSharePlugin_logic_mem_counter[8102] = 4'b0000;
    GSharePlugin_logic_mem_counter[8103] = 4'b0000;
    GSharePlugin_logic_mem_counter[8104] = 4'b0000;
    GSharePlugin_logic_mem_counter[8105] = 4'b0000;
    GSharePlugin_logic_mem_counter[8106] = 4'b0000;
    GSharePlugin_logic_mem_counter[8107] = 4'b0000;
    GSharePlugin_logic_mem_counter[8108] = 4'b0000;
    GSharePlugin_logic_mem_counter[8109] = 4'b0000;
    GSharePlugin_logic_mem_counter[8110] = 4'b0000;
    GSharePlugin_logic_mem_counter[8111] = 4'b0000;
    GSharePlugin_logic_mem_counter[8112] = 4'b0000;
    GSharePlugin_logic_mem_counter[8113] = 4'b0000;
    GSharePlugin_logic_mem_counter[8114] = 4'b0000;
    GSharePlugin_logic_mem_counter[8115] = 4'b0000;
    GSharePlugin_logic_mem_counter[8116] = 4'b0000;
    GSharePlugin_logic_mem_counter[8117] = 4'b0000;
    GSharePlugin_logic_mem_counter[8118] = 4'b0000;
    GSharePlugin_logic_mem_counter[8119] = 4'b0000;
    GSharePlugin_logic_mem_counter[8120] = 4'b0000;
    GSharePlugin_logic_mem_counter[8121] = 4'b0000;
    GSharePlugin_logic_mem_counter[8122] = 4'b0000;
    GSharePlugin_logic_mem_counter[8123] = 4'b0000;
    GSharePlugin_logic_mem_counter[8124] = 4'b0000;
    GSharePlugin_logic_mem_counter[8125] = 4'b0000;
    GSharePlugin_logic_mem_counter[8126] = 4'b0000;
    GSharePlugin_logic_mem_counter[8127] = 4'b0000;
    GSharePlugin_logic_mem_counter[8128] = 4'b0000;
    GSharePlugin_logic_mem_counter[8129] = 4'b0000;
    GSharePlugin_logic_mem_counter[8130] = 4'b0000;
    GSharePlugin_logic_mem_counter[8131] = 4'b0000;
    GSharePlugin_logic_mem_counter[8132] = 4'b0000;
    GSharePlugin_logic_mem_counter[8133] = 4'b0000;
    GSharePlugin_logic_mem_counter[8134] = 4'b0000;
    GSharePlugin_logic_mem_counter[8135] = 4'b0000;
    GSharePlugin_logic_mem_counter[8136] = 4'b0000;
    GSharePlugin_logic_mem_counter[8137] = 4'b0000;
    GSharePlugin_logic_mem_counter[8138] = 4'b0000;
    GSharePlugin_logic_mem_counter[8139] = 4'b0000;
    GSharePlugin_logic_mem_counter[8140] = 4'b0000;
    GSharePlugin_logic_mem_counter[8141] = 4'b0000;
    GSharePlugin_logic_mem_counter[8142] = 4'b0000;
    GSharePlugin_logic_mem_counter[8143] = 4'b0000;
    GSharePlugin_logic_mem_counter[8144] = 4'b0000;
    GSharePlugin_logic_mem_counter[8145] = 4'b0000;
    GSharePlugin_logic_mem_counter[8146] = 4'b0000;
    GSharePlugin_logic_mem_counter[8147] = 4'b0000;
    GSharePlugin_logic_mem_counter[8148] = 4'b0000;
    GSharePlugin_logic_mem_counter[8149] = 4'b0000;
    GSharePlugin_logic_mem_counter[8150] = 4'b0000;
    GSharePlugin_logic_mem_counter[8151] = 4'b0000;
    GSharePlugin_logic_mem_counter[8152] = 4'b0000;
    GSharePlugin_logic_mem_counter[8153] = 4'b0000;
    GSharePlugin_logic_mem_counter[8154] = 4'b0000;
    GSharePlugin_logic_mem_counter[8155] = 4'b0000;
    GSharePlugin_logic_mem_counter[8156] = 4'b0000;
    GSharePlugin_logic_mem_counter[8157] = 4'b0000;
    GSharePlugin_logic_mem_counter[8158] = 4'b0000;
    GSharePlugin_logic_mem_counter[8159] = 4'b0000;
    GSharePlugin_logic_mem_counter[8160] = 4'b0000;
    GSharePlugin_logic_mem_counter[8161] = 4'b0000;
    GSharePlugin_logic_mem_counter[8162] = 4'b0000;
    GSharePlugin_logic_mem_counter[8163] = 4'b0000;
    GSharePlugin_logic_mem_counter[8164] = 4'b0000;
    GSharePlugin_logic_mem_counter[8165] = 4'b0000;
    GSharePlugin_logic_mem_counter[8166] = 4'b0000;
    GSharePlugin_logic_mem_counter[8167] = 4'b0000;
    GSharePlugin_logic_mem_counter[8168] = 4'b0000;
    GSharePlugin_logic_mem_counter[8169] = 4'b0000;
    GSharePlugin_logic_mem_counter[8170] = 4'b0000;
    GSharePlugin_logic_mem_counter[8171] = 4'b0000;
    GSharePlugin_logic_mem_counter[8172] = 4'b0000;
    GSharePlugin_logic_mem_counter[8173] = 4'b0000;
    GSharePlugin_logic_mem_counter[8174] = 4'b0000;
    GSharePlugin_logic_mem_counter[8175] = 4'b0000;
    GSharePlugin_logic_mem_counter[8176] = 4'b0000;
    GSharePlugin_logic_mem_counter[8177] = 4'b0000;
    GSharePlugin_logic_mem_counter[8178] = 4'b0000;
    GSharePlugin_logic_mem_counter[8179] = 4'b0000;
    GSharePlugin_logic_mem_counter[8180] = 4'b0000;
    GSharePlugin_logic_mem_counter[8181] = 4'b0000;
    GSharePlugin_logic_mem_counter[8182] = 4'b0000;
    GSharePlugin_logic_mem_counter[8183] = 4'b0000;
    GSharePlugin_logic_mem_counter[8184] = 4'b0000;
    GSharePlugin_logic_mem_counter[8185] = 4'b0000;
    GSharePlugin_logic_mem_counter[8186] = 4'b0000;
    GSharePlugin_logic_mem_counter[8187] = 4'b0000;
    GSharePlugin_logic_mem_counter[8188] = 4'b0000;
    GSharePlugin_logic_mem_counter[8189] = 4'b0000;
    GSharePlugin_logic_mem_counter[8190] = 4'b0000;
    GSharePlugin_logic_mem_counter[8191] = 4'b0000;
  end
  always @(posedge clk) begin
    if(_zz_when_MultiportRam_l328) begin
      GSharePlugin_logic_mem_counter[GSharePlugin_logic_mem_write_payload_address] <= _zz_GSharePlugin_logic_mem_counter_port;
    end
  end

  always @(posedge clk) begin
    if(FetchPlugin_stages_0_ready) begin
      _zz_GSharePlugin_logic_mem_counter_port1 <= GSharePlugin_logic_mem_counter[FetchPlugin_stages_0_GSharePlugin_logic_HASH];
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_addressPre[_zz_Lsu2Plugin_logic_lq_mem_addressPre_port] <= _zz_Lsu2Plugin_logic_lq_mem_addressPre_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_addressPre_port1 = Lsu2Plugin_logic_lq_mem_addressPre[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign _zz_Lsu2Plugin_logic_lq_mem_addressPre_port2 = Lsu2Plugin_logic_lq_mem_addressPre[Lsu2Plugin_logic_lq_ptr_freeReal];
  assign _zz_Lsu2Plugin_logic_lq_mem_addressPost_port0 = Lsu2Plugin_logic_lq_mem_addressPost[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(_zz_13) begin
      Lsu2Plugin_logic_lq_mem_addressPost[Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID] <= _zz_Lsu2Plugin_logic_lq_mem_addressPost_port;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_addressPost_port2 = Lsu2Plugin_logic_lq_mem_addressPost[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_size[_zz_Lsu2Plugin_logic_lq_mem_size_port] <= _zz_Lsu2Plugin_logic_lq_mem_size_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_size_port1 = Lsu2Plugin_logic_lq_mem_size[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign _zz_Lsu2Plugin_logic_lq_mem_size_port2 = Lsu2Plugin_logic_lq_mem_size[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_physRd[_zz_Lsu2Plugin_logic_lq_mem_physRd_port] <= _zz_Lsu2Plugin_logic_lq_mem_physRd_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_physRd_port1 = Lsu2Plugin_logic_lq_mem_physRd[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign _zz_Lsu2Plugin_logic_lq_mem_physRd_port2 = Lsu2Plugin_logic_lq_mem_physRd[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_robId[_zz_Lsu2Plugin_logic_lq_mem_robId_port] <= _zz_Lsu2Plugin_logic_lq_mem_robId_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_robId_port1 = Lsu2Plugin_logic_lq_mem_robId[Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID];
  assign _zz_Lsu2Plugin_logic_lq_mem_robId_port2 = Lsu2Plugin_logic_lq_mem_robId[Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel];
  assign _zz_Lsu2Plugin_logic_lq_mem_robId_port3 = Lsu2Plugin_logic_lq_mem_robId[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_robIdMsb[_zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port] <= _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port1 = Lsu2Plugin_logic_lq_mem_robIdMsb[Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_pc[_zz_Lsu2Plugin_logic_lq_mem_pc_port] <= _zz_Lsu2Plugin_logic_lq_mem_pc_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_pc_port1 = Lsu2Plugin_logic_lq_mem_pc[_zz_Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC];
  assign _zz_Lsu2Plugin_logic_lq_mem_io_port0 = Lsu2Plugin_logic_lq_mem_io[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(_zz_12) begin
      Lsu2Plugin_logic_lq_mem_io[Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID] <= _zz_Lsu2Plugin_logic_lq_mem_io_port;
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_writeRd[_zz_Lsu2Plugin_logic_lq_mem_writeRd_port] <= _zz_Lsu2Plugin_logic_lq_mem_writeRd_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_writeRd_port1 = Lsu2Plugin_logic_lq_mem_writeRd[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign _zz_Lsu2Plugin_logic_lq_mem_writeRd_port2 = Lsu2Plugin_logic_lq_mem_writeRd[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_lr[_zz_Lsu2Plugin_logic_lq_mem_lr_port] <= _zz_Lsu2Plugin_logic_lq_mem_lr_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_lr_port1 = Lsu2Plugin_logic_lq_mem_lr[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_unsigned[_zz_Lsu2Plugin_logic_lq_mem_unsigned_port] <= _zz_Lsu2Plugin_logic_lq_mem_unsigned_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_unsigned_port1 = Lsu2Plugin_logic_lq_mem_unsigned[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  assign _zz_Lsu2Plugin_logic_lq_mem_unsigned_port2 = Lsu2Plugin_logic_lq_mem_unsigned[Lsu2Plugin_logic_lq_ptr_freeReal];
  always @(posedge clk) begin
    if(_zz_15) begin
      Lsu2Plugin_logic_lq_mem_spFpAddress[FrontendPlugin_dispatch_LQ_ID_0] <= _zz_Lsu2Plugin_logic_lq_mem_spFpAddress_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_14) begin
      Lsu2Plugin_logic_lq_mem_spFpAddress[FrontendPlugin_dispatch_LQ_ID_1] <= _zz_Lsu2Plugin_logic_lq_mem_spFpAddress_port_1;
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_hazardPrediction_valid[_zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port] <= _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port1 = Lsu2Plugin_logic_lq_mem_hazardPrediction_valid[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_hazardPrediction_delta[_zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port] <= _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port1 = Lsu2Plugin_logic_lq_mem_hazardPrediction_delta[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_hazardPrediction_score[_zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port] <= _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port1 = Lsu2Plugin_logic_lq_mem_hazardPrediction_score[Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      Lsu2Plugin_logic_lq_mem_hitPrediction_counter[_zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port] <= _zz_Lsu2Plugin_logic_lq_mem_hitPrediction_counter_port_1;
    end
  end

  initial begin
    Lsu2Plugin_logic_lq_hazardPrediction_mem[0] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[1] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[2] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[3] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[4] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[5] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[6] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[7] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[8] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[9] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[10] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[11] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[12] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[13] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[14] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[15] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[16] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[17] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[18] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[19] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[20] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[21] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[22] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[23] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[24] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[25] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[26] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[27] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[28] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[29] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[30] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[31] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[32] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[33] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[34] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[35] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[36] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[37] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[38] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[39] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[40] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[41] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[42] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[43] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[44] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[45] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[46] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[47] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[48] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[49] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[50] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[51] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[52] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[53] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[54] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[55] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[56] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[57] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[58] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[59] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[60] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[61] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[62] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[63] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[64] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[65] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[66] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[67] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[68] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[69] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[70] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[71] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[72] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[73] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[74] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[75] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[76] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[77] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[78] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[79] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[80] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[81] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[82] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[83] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[84] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[85] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[86] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[87] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[88] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[89] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[90] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[91] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[92] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[93] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[94] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[95] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[96] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[97] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[98] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[99] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[100] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[101] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[102] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[103] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[104] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[105] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[106] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[107] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[108] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[109] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[110] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[111] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[112] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[113] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[114] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[115] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[116] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[117] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[118] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[119] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[120] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[121] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[122] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[123] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[124] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[125] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[126] = 23'b00000000000000000000000;
    Lsu2Plugin_logic_lq_hazardPrediction_mem[127] = 23'b00000000000000000000000;
  end
  always @(posedge clk) begin
    if(_zz_when_MultiportRam_l362_1) begin
      Lsu2Plugin_logic_lq_hazardPrediction_mem[_zz_when_MultiportRam_l362_2] <= _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_valid) begin
      _zz_Lsu2Plugin_logic_lq_hazardPrediction_mem_port1 <= Lsu2Plugin_logic_lq_hazardPrediction_mem[Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_payload];
    end
  end

  initial begin
    Lsu2Plugin_logic_lq_hitPrediction_mem[0] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[2] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[3] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[4] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[5] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[6] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[7] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[8] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[9] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[10] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[11] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[12] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[13] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[14] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[15] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[16] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[17] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[18] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[19] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[20] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[21] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[22] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[23] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[24] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[25] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[26] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[27] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[28] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[29] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[30] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[31] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[32] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[33] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[34] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[35] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[36] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[37] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[38] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[39] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[40] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[41] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[42] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[43] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[44] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[45] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[46] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[47] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[48] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[49] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[50] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[51] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[52] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[53] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[54] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[55] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[56] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[57] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[58] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[59] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[60] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[61] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[62] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[63] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[64] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[65] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[66] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[67] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[68] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[69] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[70] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[71] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[72] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[73] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[74] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[75] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[76] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[77] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[78] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[79] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[80] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[81] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[82] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[83] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[84] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[85] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[86] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[87] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[88] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[89] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[90] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[91] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[92] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[93] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[94] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[95] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[96] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[97] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[98] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[99] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[100] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[101] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[102] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[103] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[104] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[105] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[106] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[107] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[108] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[109] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[110] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[111] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[112] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[113] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[114] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[115] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[116] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[117] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[118] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[119] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[120] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[121] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[122] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[123] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[124] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[125] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[126] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[127] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[128] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[129] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[130] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[131] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[132] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[133] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[134] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[135] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[136] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[137] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[138] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[139] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[140] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[141] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[142] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[143] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[144] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[145] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[146] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[147] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[148] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[149] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[150] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[151] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[152] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[153] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[154] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[155] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[156] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[157] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[158] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[159] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[160] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[161] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[162] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[163] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[164] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[165] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[166] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[167] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[168] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[169] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[170] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[171] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[172] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[173] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[174] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[175] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[176] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[177] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[178] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[179] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[180] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[181] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[182] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[183] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[184] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[185] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[186] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[187] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[188] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[189] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[190] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[191] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[192] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[193] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[194] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[195] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[196] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[197] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[198] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[199] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[200] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[201] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[202] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[203] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[204] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[205] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[206] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[207] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[208] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[209] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[210] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[211] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[212] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[213] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[214] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[215] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[216] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[217] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[218] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[219] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[220] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[221] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[222] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[223] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[224] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[225] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[226] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[227] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[228] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[229] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[230] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[231] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[232] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[233] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[234] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[235] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[236] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[237] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[238] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[239] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[240] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[241] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[242] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[243] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[244] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[245] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[246] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[247] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[248] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[249] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[250] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[251] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[252] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[253] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[254] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[255] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[256] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[257] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[258] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[259] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[260] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[261] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[262] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[263] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[264] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[265] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[266] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[267] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[268] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[269] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[270] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[271] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[272] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[273] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[274] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[275] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[276] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[277] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[278] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[279] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[280] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[281] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[282] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[283] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[284] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[285] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[286] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[287] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[288] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[289] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[290] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[291] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[292] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[293] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[294] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[295] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[296] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[297] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[298] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[299] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[300] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[301] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[302] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[303] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[304] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[305] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[306] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[307] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[308] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[309] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[310] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[311] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[312] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[313] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[314] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[315] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[316] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[317] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[318] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[319] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[320] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[321] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[322] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[323] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[324] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[325] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[326] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[327] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[328] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[329] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[330] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[331] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[332] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[333] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[334] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[335] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[336] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[337] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[338] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[339] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[340] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[341] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[342] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[343] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[344] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[345] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[346] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[347] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[348] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[349] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[350] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[351] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[352] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[353] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[354] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[355] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[356] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[357] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[358] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[359] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[360] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[361] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[362] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[363] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[364] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[365] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[366] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[367] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[368] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[369] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[370] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[371] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[372] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[373] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[374] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[375] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[376] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[377] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[378] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[379] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[380] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[381] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[382] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[383] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[384] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[385] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[386] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[387] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[388] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[389] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[390] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[391] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[392] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[393] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[394] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[395] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[396] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[397] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[398] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[399] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[400] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[401] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[402] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[403] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[404] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[405] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[406] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[407] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[408] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[409] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[410] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[411] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[412] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[413] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[414] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[415] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[416] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[417] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[418] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[419] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[420] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[421] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[422] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[423] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[424] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[425] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[426] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[427] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[428] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[429] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[430] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[431] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[432] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[433] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[434] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[435] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[436] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[437] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[438] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[439] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[440] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[441] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[442] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[443] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[444] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[445] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[446] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[447] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[448] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[449] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[450] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[451] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[452] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[453] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[454] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[455] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[456] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[457] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[458] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[459] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[460] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[461] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[462] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[463] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[464] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[465] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[466] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[467] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[468] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[469] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[470] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[471] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[472] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[473] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[474] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[475] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[476] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[477] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[478] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[479] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[480] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[481] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[482] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[483] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[484] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[485] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[486] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[487] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[488] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[489] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[490] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[491] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[492] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[493] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[494] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[495] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[496] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[497] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[498] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[499] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[500] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[501] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[502] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[503] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[504] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[505] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[506] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[507] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[508] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[509] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[510] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[511] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[512] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[513] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[514] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[515] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[516] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[517] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[518] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[519] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[520] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[521] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[522] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[523] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[524] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[525] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[526] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[527] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[528] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[529] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[530] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[531] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[532] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[533] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[534] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[535] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[536] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[537] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[538] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[539] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[540] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[541] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[542] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[543] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[544] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[545] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[546] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[547] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[548] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[549] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[550] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[551] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[552] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[553] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[554] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[555] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[556] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[557] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[558] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[559] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[560] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[561] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[562] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[563] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[564] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[565] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[566] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[567] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[568] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[569] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[570] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[571] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[572] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[573] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[574] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[575] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[576] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[577] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[578] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[579] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[580] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[581] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[582] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[583] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[584] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[585] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[586] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[587] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[588] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[589] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[590] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[591] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[592] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[593] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[594] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[595] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[596] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[597] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[598] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[599] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[600] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[601] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[602] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[603] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[604] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[605] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[606] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[607] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[608] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[609] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[610] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[611] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[612] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[613] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[614] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[615] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[616] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[617] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[618] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[619] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[620] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[621] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[622] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[623] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[624] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[625] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[626] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[627] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[628] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[629] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[630] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[631] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[632] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[633] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[634] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[635] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[636] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[637] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[638] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[639] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[640] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[641] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[642] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[643] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[644] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[645] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[646] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[647] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[648] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[649] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[650] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[651] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[652] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[653] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[654] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[655] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[656] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[657] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[658] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[659] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[660] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[661] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[662] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[663] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[664] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[665] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[666] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[667] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[668] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[669] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[670] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[671] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[672] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[673] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[674] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[675] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[676] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[677] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[678] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[679] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[680] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[681] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[682] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[683] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[684] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[685] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[686] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[687] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[688] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[689] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[690] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[691] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[692] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[693] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[694] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[695] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[696] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[697] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[698] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[699] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[700] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[701] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[702] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[703] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[704] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[705] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[706] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[707] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[708] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[709] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[710] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[711] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[712] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[713] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[714] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[715] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[716] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[717] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[718] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[719] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[720] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[721] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[722] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[723] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[724] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[725] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[726] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[727] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[728] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[729] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[730] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[731] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[732] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[733] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[734] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[735] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[736] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[737] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[738] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[739] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[740] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[741] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[742] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[743] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[744] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[745] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[746] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[747] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[748] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[749] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[750] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[751] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[752] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[753] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[754] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[755] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[756] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[757] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[758] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[759] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[760] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[761] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[762] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[763] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[764] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[765] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[766] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[767] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[768] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[769] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[770] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[771] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[772] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[773] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[774] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[775] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[776] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[777] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[778] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[779] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[780] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[781] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[782] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[783] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[784] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[785] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[786] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[787] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[788] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[789] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[790] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[791] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[792] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[793] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[794] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[795] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[796] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[797] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[798] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[799] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[800] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[801] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[802] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[803] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[804] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[805] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[806] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[807] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[808] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[809] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[810] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[811] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[812] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[813] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[814] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[815] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[816] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[817] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[818] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[819] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[820] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[821] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[822] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[823] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[824] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[825] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[826] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[827] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[828] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[829] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[830] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[831] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[832] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[833] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[834] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[835] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[836] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[837] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[838] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[839] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[840] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[841] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[842] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[843] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[844] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[845] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[846] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[847] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[848] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[849] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[850] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[851] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[852] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[853] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[854] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[855] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[856] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[857] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[858] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[859] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[860] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[861] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[862] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[863] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[864] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[865] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[866] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[867] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[868] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[869] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[870] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[871] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[872] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[873] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[874] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[875] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[876] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[877] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[878] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[879] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[880] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[881] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[882] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[883] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[884] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[885] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[886] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[887] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[888] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[889] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[890] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[891] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[892] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[893] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[894] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[895] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[896] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[897] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[898] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[899] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[900] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[901] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[902] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[903] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[904] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[905] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[906] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[907] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[908] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[909] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[910] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[911] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[912] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[913] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[914] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[915] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[916] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[917] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[918] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[919] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[920] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[921] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[922] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[923] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[924] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[925] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[926] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[927] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[928] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[929] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[930] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[931] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[932] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[933] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[934] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[935] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[936] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[937] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[938] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[939] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[940] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[941] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[942] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[943] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[944] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[945] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[946] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[947] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[948] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[949] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[950] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[951] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[952] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[953] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[954] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[955] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[956] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[957] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[958] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[959] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[960] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[961] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[962] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[963] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[964] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[965] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[966] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[967] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[968] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[969] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[970] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[971] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[972] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[973] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[974] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[975] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[976] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[977] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[978] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[979] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[980] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[981] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[982] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[983] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[984] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[985] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[986] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[987] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[988] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[989] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[990] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[991] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[992] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[993] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[994] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[995] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[996] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[997] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[998] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[999] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1000] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1001] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1002] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1003] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1004] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1005] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1006] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1007] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1008] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1009] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1010] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1011] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1012] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1013] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1014] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1015] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1016] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1017] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1018] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1019] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1020] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1021] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1022] = 6'b000000;
    Lsu2Plugin_logic_lq_hitPrediction_mem[1023] = 6'b000000;
  end
  always @(posedge clk) begin
    if(_zz_when_MultiportRam_l362) begin
      Lsu2Plugin_logic_lq_hitPrediction_mem[_zz_when_MultiportRam_l362_3] <= _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter;
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_valid) begin
      _zz_Lsu2Plugin_logic_lq_hitPrediction_mem_port1 <= Lsu2Plugin_logic_lq_hitPrediction_mem[Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_robId[_zz_Lsu2Plugin_logic_sq_mem_robId_port] <= _zz_Lsu2Plugin_logic_sq_mem_robId_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_robId_port1 = Lsu2Plugin_logic_sq_mem_robId[Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID];
  assign _zz_Lsu2Plugin_logic_sq_mem_robId_port2 = Lsu2Plugin_logic_sq_mem_robId[Lsu2Plugin_logic_sq_ptr_commitReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_robIdMsb[_zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port] <= _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port1 = Lsu2Plugin_logic_sq_mem_robIdMsb[Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_addressPre[_zz_Lsu2Plugin_logic_sq_mem_addressPre_port] <= _zz_Lsu2Plugin_logic_sq_mem_addressPre_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_addressPre_port1 = Lsu2Plugin_logic_sq_mem_addressPre[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  assign _zz_Lsu2Plugin_logic_sq_mem_addressPre_port2 = Lsu2Plugin_logic_sq_mem_addressPre[Lsu2Plugin_logic_sq_ptr_commitReal];
  assign _zz_Lsu2Plugin_logic_sq_mem_addressPost_port0 = Lsu2Plugin_logic_sq_mem_addressPost[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  always @(posedge clk) begin
    if(_zz_11) begin
      Lsu2Plugin_logic_sq_mem_addressPost[Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID] <= _zz_Lsu2Plugin_logic_sq_mem_addressPost_port;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_addressPost_port2 = Lsu2Plugin_logic_sq_mem_addressPost[Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID];
  assign _zz_Lsu2Plugin_logic_sq_mem_addressPost_port3 = Lsu2Plugin_logic_sq_mem_addressPost[Lsu2Plugin_logic_sq_ptr_writeBackReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_size[_zz_Lsu2Plugin_logic_sq_mem_size_port] <= _zz_Lsu2Plugin_logic_sq_mem_size_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_size_port1 = Lsu2Plugin_logic_sq_mem_size[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  assign _zz_Lsu2Plugin_logic_sq_mem_size_port2 = Lsu2Plugin_logic_sq_mem_size[Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID];
  assign _zz_Lsu2Plugin_logic_sq_mem_size_port3 = Lsu2Plugin_logic_sq_mem_size[Lsu2Plugin_logic_sq_ptr_writeBackReal];
  assign _zz_Lsu2Plugin_logic_sq_mem_size_port4 = Lsu2Plugin_logic_sq_mem_size[Lsu2Plugin_logic_sq_ptr_commitReal];
  assign _zz_Lsu2Plugin_logic_sq_mem_io_port0 = Lsu2Plugin_logic_sq_mem_io[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  always @(posedge clk) begin
    if(_zz_10) begin
      Lsu2Plugin_logic_sq_mem_io[Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID] <= _zz_Lsu2Plugin_logic_sq_mem_io_port;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_io_port2 = Lsu2Plugin_logic_sq_mem_io[Lsu2Plugin_logic_sq_ptr_writeBackReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_amo[_zz_Lsu2Plugin_logic_sq_mem_amo_port] <= _zz_Lsu2Plugin_logic_sq_mem_amo_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_amo_port1 = Lsu2Plugin_logic_sq_mem_amo[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  assign _zz_Lsu2Plugin_logic_sq_mem_amo_port2 = Lsu2Plugin_logic_sq_mem_amo[Lsu2Plugin_logic_sq_ptr_commitReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_sc[_zz_Lsu2Plugin_logic_sq_mem_sc_port] <= _zz_Lsu2Plugin_logic_sq_mem_sc_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_sc_port1 = Lsu2Plugin_logic_sq_mem_sc[Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID];
  assign _zz_Lsu2Plugin_logic_sq_mem_sc_port2 = Lsu2Plugin_logic_sq_mem_sc[Lsu2Plugin_logic_sq_ptr_commitReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_data[_zz_Lsu2Plugin_logic_sq_mem_data_port] <= AguPlugin_setup_port_payload_data;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_data_port1 = Lsu2Plugin_logic_sq_mem_data[Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID];
  assign _zz_Lsu2Plugin_logic_sq_mem_data_port2 = Lsu2Plugin_logic_sq_mem_data[Lsu2Plugin_logic_sq_ptr_writeBackReal];
  always @(posedge clk) begin
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      Lsu2Plugin_logic_sq_mem_doNotBypass[_zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port] <= _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port_1;
    end
  end

  assign _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port1 = Lsu2Plugin_logic_sq_mem_doNotBypass[Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0[FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port;
    end
  end

  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0[FetchCachePlugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1[FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port;
    end
  end

  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1[FetchCachePlugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2[FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port;
    end
  end

  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2[FetchCachePlugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3[FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port;
    end
  end

  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3[FetchCachePlugin_logic_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0[FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port;
    end
  end

  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0[FetchCachePlugin_logic_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port_1) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1[FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address] <= _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port;
    end
  end

  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port1 = FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1[FetchCachePlugin_logic_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0[Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port;
    end
  end

  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1[Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port;
    end
  end

  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2[Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port;
    end
  end

  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3[Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port;
    end
  end

  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0[Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port;
    end
  end

  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port_1) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1[Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address] <= _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port;
    end
  end

  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port1 = Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1[Lsu2Plugin_logic_sharedPip_translationPort_logic_read_1_readAddress];
  always @(posedge clk) begin
    if(_zz_9) begin
      CsrRamPlugin_logic_mem[CsrRamPlugin_logic_writeLogic_port_payload_address] <= CsrRamPlugin_logic_writeLogic_port_payload_data;
    end
  end

  assign _zz_CsrRamPlugin_logic_mem_port1 = CsrRamPlugin_logic_mem[CsrRamPlugin_logic_readLogic_port_address];
  always @(posedge clk) begin
    if(_zz_8) begin
      RobPlugin_logic_completionMem_target[RobPlugin_logic_completionMem_targetWrite_payload_address] <= RobPlugin_logic_completionMem_targetWrite_payload_data;
    end
  end

  assign _zz_RobPlugin_logic_completionMem_target_port1 = RobPlugin_logic_completionMem_target[RobPlugin_logic_completionMem_reads_0_targetRead_address];
  initial begin
    RobPlugin_logic_completionMem_hits_0[0] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[1] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[2] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[3] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[4] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[5] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[6] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[7] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[8] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[9] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[10] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[11] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[12] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[13] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[14] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[15] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[16] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[17] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[18] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[19] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[20] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[21] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[22] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[23] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[24] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[25] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[26] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[27] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[28] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[29] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[30] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[31] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[32] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[33] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[34] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[35] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[36] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[37] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[38] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[39] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[40] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[41] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[42] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[43] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[44] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[45] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[46] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[47] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[48] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[49] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[50] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[51] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[52] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[53] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[54] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[55] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[56] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[57] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[58] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[59] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[60] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[61] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[62] = 1'b0;
    RobPlugin_logic_completionMem_hits_0[63] = 1'b0;
  end
  assign _zz_RobPlugin_logic_completionMem_hits_0_port0 = RobPlugin_logic_completionMem_hits_0[RobPlugin_logic_completionMem_init_0_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_0_port1 = RobPlugin_logic_completionMem_hits_0[RobPlugin_logic_completionMem_init_1_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_0_port2 = RobPlugin_logic_completionMem_hits_0[Lsu2Plugin_setup_sharedCompletion_payload_id];
  always @(posedge clk) begin
    if(_zz_7) begin
      RobPlugin_logic_completionMem_hits_0[Lsu2Plugin_setup_sharedCompletion_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_0_port;
    end
  end

  assign _zz_RobPlugin_logic_completionMem_hits_0_port4 = RobPlugin_logic_completionMem_hits_0[_zz_CommitPlugin_setup_robLineMask_mask];
  assign _zz_RobPlugin_logic_completionMem_hits_0_port5 = RobPlugin_logic_completionMem_hits_0[_zz_CommitPlugin_setup_robLineMask_mask_1];
  initial begin
    RobPlugin_logic_completionMem_hits_1[0] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[1] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[2] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[3] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[4] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[5] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[6] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[7] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[8] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[9] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[10] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[11] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[12] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[13] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[14] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[15] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[16] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[17] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[18] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[19] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[20] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[21] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[22] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[23] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[24] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[25] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[26] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[27] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[28] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[29] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[30] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[31] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[32] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[33] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[34] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[35] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[36] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[37] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[38] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[39] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[40] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[41] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[42] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[43] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[44] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[45] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[46] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[47] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[48] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[49] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[50] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[51] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[52] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[53] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[54] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[55] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[56] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[57] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[58] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[59] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[60] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[61] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[62] = 1'b0;
    RobPlugin_logic_completionMem_hits_1[63] = 1'b0;
  end
  assign _zz_RobPlugin_logic_completionMem_hits_1_port0 = RobPlugin_logic_completionMem_hits_1[RobPlugin_logic_completionMem_init_0_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_1_port1 = RobPlugin_logic_completionMem_hits_1[RobPlugin_logic_completionMem_init_1_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_1_port2 = RobPlugin_logic_completionMem_hits_1[Lsu2Plugin_setup_specialCompletion_payload_id];
  always @(posedge clk) begin
    if(_zz_6) begin
      RobPlugin_logic_completionMem_hits_1[Lsu2Plugin_setup_specialCompletion_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_1_port;
    end
  end

  assign _zz_RobPlugin_logic_completionMem_hits_1_port4 = RobPlugin_logic_completionMem_hits_1[_zz_CommitPlugin_setup_robLineMask_mask];
  assign _zz_RobPlugin_logic_completionMem_hits_1_port5 = RobPlugin_logic_completionMem_hits_1[_zz_CommitPlugin_setup_robLineMask_mask_1];
  initial begin
    RobPlugin_logic_completionMem_hits_2[0] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[1] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[2] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[3] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[4] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[5] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[6] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[7] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[8] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[9] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[10] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[11] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[12] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[13] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[14] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[15] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[16] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[17] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[18] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[19] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[20] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[21] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[22] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[23] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[24] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[25] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[26] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[27] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[28] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[29] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[30] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[31] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[32] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[33] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[34] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[35] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[36] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[37] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[38] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[39] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[40] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[41] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[42] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[43] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[44] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[45] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[46] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[47] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[48] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[49] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[50] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[51] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[52] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[53] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[54] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[55] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[56] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[57] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[58] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[59] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[60] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[61] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[62] = 1'b0;
    RobPlugin_logic_completionMem_hits_2[63] = 1'b0;
  end
  assign _zz_RobPlugin_logic_completionMem_hits_2_port0 = RobPlugin_logic_completionMem_hits_2[RobPlugin_logic_completionMem_init_0_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_2_port1 = RobPlugin_logic_completionMem_hits_2[RobPlugin_logic_completionMem_init_1_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_2_port2 = RobPlugin_logic_completionMem_hits_2[ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id];
  always @(posedge clk) begin
    if(_zz_5) begin
      RobPlugin_logic_completionMem_hits_2[ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_2_port;
    end
  end

  assign _zz_RobPlugin_logic_completionMem_hits_2_port4 = RobPlugin_logic_completionMem_hits_2[_zz_CommitPlugin_setup_robLineMask_mask];
  assign _zz_RobPlugin_logic_completionMem_hits_2_port5 = RobPlugin_logic_completionMem_hits_2[_zz_CommitPlugin_setup_robLineMask_mask_1];
  initial begin
    RobPlugin_logic_completionMem_hits_3[0] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[1] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[2] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[3] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[4] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[5] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[6] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[7] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[8] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[9] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[10] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[11] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[12] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[13] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[14] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[15] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[16] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[17] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[18] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[19] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[20] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[21] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[22] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[23] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[24] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[25] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[26] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[27] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[28] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[29] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[30] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[31] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[32] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[33] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[34] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[35] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[36] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[37] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[38] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[39] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[40] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[41] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[42] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[43] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[44] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[45] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[46] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[47] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[48] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[49] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[50] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[51] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[52] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[53] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[54] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[55] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[56] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[57] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[58] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[59] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[60] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[61] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[62] = 1'b0;
    RobPlugin_logic_completionMem_hits_3[63] = 1'b0;
  end
  assign _zz_RobPlugin_logic_completionMem_hits_3_port0 = RobPlugin_logic_completionMem_hits_3[RobPlugin_logic_completionMem_init_0_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_3_port1 = RobPlugin_logic_completionMem_hits_3[RobPlugin_logic_completionMem_init_1_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_3_port2 = RobPlugin_logic_completionMem_hits_3[ALU0_ExecutionUnitBase_pipeline_completion_1_port_payload_id];
  always @(posedge clk) begin
    if(_zz_4) begin
      RobPlugin_logic_completionMem_hits_3[ALU0_ExecutionUnitBase_pipeline_completion_1_port_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_3_port;
    end
  end

  assign _zz_RobPlugin_logic_completionMem_hits_3_port4 = RobPlugin_logic_completionMem_hits_3[_zz_CommitPlugin_setup_robLineMask_mask];
  assign _zz_RobPlugin_logic_completionMem_hits_3_port5 = RobPlugin_logic_completionMem_hits_3[_zz_CommitPlugin_setup_robLineMask_mask_1];
  initial begin
    RobPlugin_logic_completionMem_hits_4[0] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[1] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[2] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[3] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[4] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[5] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[6] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[7] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[8] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[9] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[10] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[11] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[12] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[13] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[14] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[15] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[16] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[17] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[18] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[19] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[20] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[21] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[22] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[23] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[24] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[25] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[26] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[27] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[28] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[29] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[30] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[31] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[32] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[33] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[34] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[35] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[36] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[37] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[38] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[39] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[40] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[41] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[42] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[43] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[44] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[45] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[46] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[47] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[48] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[49] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[50] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[51] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[52] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[53] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[54] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[55] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[56] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[57] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[58] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[59] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[60] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[61] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[62] = 1'b0;
    RobPlugin_logic_completionMem_hits_4[63] = 1'b0;
  end
  assign _zz_RobPlugin_logic_completionMem_hits_4_port0 = RobPlugin_logic_completionMem_hits_4[RobPlugin_logic_completionMem_init_0_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_4_port1 = RobPlugin_logic_completionMem_hits_4[RobPlugin_logic_completionMem_init_1_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_4_port2 = RobPlugin_logic_completionMem_hits_4[ALU1_ExecutionUnitBase_pipeline_completion_0_port_payload_id];
  always @(posedge clk) begin
    if(_zz_3) begin
      RobPlugin_logic_completionMem_hits_4[ALU1_ExecutionUnitBase_pipeline_completion_0_port_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_4_port;
    end
  end

  assign _zz_RobPlugin_logic_completionMem_hits_4_port4 = RobPlugin_logic_completionMem_hits_4[_zz_CommitPlugin_setup_robLineMask_mask];
  assign _zz_RobPlugin_logic_completionMem_hits_4_port5 = RobPlugin_logic_completionMem_hits_4[_zz_CommitPlugin_setup_robLineMask_mask_1];
  initial begin
    RobPlugin_logic_completionMem_hits_5[0] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[1] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[2] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[3] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[4] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[5] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[6] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[7] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[8] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[9] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[10] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[11] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[12] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[13] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[14] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[15] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[16] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[17] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[18] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[19] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[20] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[21] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[22] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[23] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[24] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[25] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[26] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[27] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[28] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[29] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[30] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[31] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[32] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[33] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[34] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[35] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[36] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[37] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[38] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[39] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[40] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[41] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[42] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[43] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[44] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[45] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[46] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[47] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[48] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[49] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[50] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[51] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[52] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[53] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[54] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[55] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[56] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[57] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[58] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[59] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[60] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[61] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[62] = 1'b0;
    RobPlugin_logic_completionMem_hits_5[63] = 1'b0;
  end
  assign _zz_RobPlugin_logic_completionMem_hits_5_port0 = RobPlugin_logic_completionMem_hits_5[RobPlugin_logic_completionMem_init_0_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_5_port1 = RobPlugin_logic_completionMem_hits_5[RobPlugin_logic_completionMem_init_1_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_5_port2 = RobPlugin_logic_completionMem_hits_5[ALU1_ExecutionUnitBase_pipeline_completion_1_port_payload_id];
  always @(posedge clk) begin
    if(_zz_2) begin
      RobPlugin_logic_completionMem_hits_5[ALU1_ExecutionUnitBase_pipeline_completion_1_port_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_5_port;
    end
  end

  assign _zz_RobPlugin_logic_completionMem_hits_5_port4 = RobPlugin_logic_completionMem_hits_5[_zz_CommitPlugin_setup_robLineMask_mask];
  assign _zz_RobPlugin_logic_completionMem_hits_5_port5 = RobPlugin_logic_completionMem_hits_5[_zz_CommitPlugin_setup_robLineMask_mask_1];
  initial begin
    RobPlugin_logic_completionMem_hits_6[0] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[1] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[2] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[3] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[4] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[5] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[6] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[7] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[8] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[9] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[10] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[11] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[12] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[13] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[14] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[15] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[16] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[17] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[18] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[19] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[20] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[21] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[22] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[23] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[24] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[25] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[26] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[27] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[28] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[29] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[30] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[31] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[32] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[33] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[34] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[35] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[36] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[37] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[38] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[39] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[40] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[41] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[42] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[43] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[44] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[45] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[46] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[47] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[48] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[49] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[50] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[51] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[52] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[53] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[54] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[55] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[56] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[57] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[58] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[59] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[60] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[61] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[62] = 1'b0;
    RobPlugin_logic_completionMem_hits_6[63] = 1'b0;
  end
  assign _zz_RobPlugin_logic_completionMem_hits_6_port0 = RobPlugin_logic_completionMem_hits_6[RobPlugin_logic_completionMem_init_0_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_6_port1 = RobPlugin_logic_completionMem_hits_6[RobPlugin_logic_completionMem_init_1_robId];
  assign _zz_RobPlugin_logic_completionMem_hits_6_port2 = RobPlugin_logic_completionMem_hits_6[EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id];
  always @(posedge clk) begin
    if(_zz_1) begin
      RobPlugin_logic_completionMem_hits_6[EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id] <= _zz_RobPlugin_logic_completionMem_hits_6_port;
    end
  end

  assign _zz_RobPlugin_logic_completionMem_hits_6_port4 = RobPlugin_logic_completionMem_hits_6[_zz_CommitPlugin_setup_robLineMask_mask];
  assign _zz_RobPlugin_logic_completionMem_hits_6_port5 = RobPlugin_logic_completionMem_hits_6[_zz_CommitPlugin_setup_robLineMask_mask_1];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port_2) begin
      RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0[_zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port] <= _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port_1;
    end
  end

  assign _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port1 = RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0[_zz_CommitPlugin_logic_commit_active];
  assign _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port2 = RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0[_zz_integer_RfAllocationPlugin_logic_push_mask_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PC_banks_0_port_1) begin
      RobPlugin_logic_storage_PC_banks_0[_zz_224] <= _zz_RobPlugin_logic_storage_PC_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_PC_banks_0_port1 = RobPlugin_logic_storage_PC_banks_0[_zz_commit_pc_0];
  assign _zz_RobPlugin_logic_storage_PC_banks_0_port2 = RobPlugin_logic_storage_PC_banks_0[_zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc];
  assign _zz_RobPlugin_logic_storage_PC_banks_0_port3 = RobPlugin_logic_storage_PC_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC];
  assign _zz_RobPlugin_logic_storage_PC_banks_0_port4 = RobPlugin_logic_storage_PC_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PC_banks_1_port_1) begin
      RobPlugin_logic_storage_PC_banks_1[_zz_224] <= _zz_RobPlugin_logic_storage_PC_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_PC_banks_1_port1 = RobPlugin_logic_storage_PC_banks_1[_zz_commit_pc_0];
  assign _zz_RobPlugin_logic_storage_PC_banks_1_port2 = RobPlugin_logic_storage_PC_banks_1[_zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc];
  assign _zz_RobPlugin_logic_storage_PC_banks_1_port3 = RobPlugin_logic_storage_PC_banks_1[_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PC];
  assign _zz_RobPlugin_logic_storage_PC_banks_1_port4 = RobPlugin_logic_storage_PC_banks_1[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port_1) begin
      RobPlugin_logic_storage_WRITE_RD_banks_0[_zz_235] <= _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port1 = RobPlugin_logic_storage_WRITE_RD_banks_0[_zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0];
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port2 = RobPlugin_logic_storage_WRITE_RD_banks_0[_zz_integer_RfAllocationPlugin_logic_push_writeRd_0];
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port3 = RobPlugin_logic_storage_WRITE_RD_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD];
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port4 = RobPlugin_logic_storage_WRITE_RD_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port_1) begin
      RobPlugin_logic_storage_WRITE_RD_banks_1[_zz_235] <= _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port1 = RobPlugin_logic_storage_WRITE_RD_banks_1[_zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0];
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port2 = RobPlugin_logic_storage_WRITE_RD_banks_1[_zz_integer_RfAllocationPlugin_logic_push_writeRd_0];
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port3 = RobPlugin_logic_storage_WRITE_RD_banks_1[_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD];
  assign _zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port4 = RobPlugin_logic_storage_WRITE_RD_banks_1[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port_2) begin
      RobPlugin_logic_storage_PHYS_RD_banks_0[_zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port] <= _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port_1;
    end
  end

  assign _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port1 = RobPlugin_logic_storage_PHYS_RD_banks_0[_zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0];
  assign _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port2 = RobPlugin_logic_storage_PHYS_RD_banks_0[_zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port_2) begin
      RobPlugin_logic_storage_ARCH_RD_banks_0[_zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port] <= _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port_1;
    end
  end

  assign _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port1 = RobPlugin_logic_storage_ARCH_RD_banks_0[_zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port_2) begin
      RobPlugin_logic_storage_PHYS_RD_FREE_banks_0[_zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port] <= _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port_1;
    end
  end

  assign _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port1 = RobPlugin_logic_storage_PHYS_RD_FREE_banks_0[_zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port_2) begin
      RobPlugin_logic_storage_BRANCH_SEL_banks_0[_zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port] <= _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port_1;
    end
  end

  assign _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port1 = RobPlugin_logic_storage_BRANCH_SEL_banks_0[_zz_BranchContextPlugin_logic_onCommit_isBranch_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port_1) begin
      RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0[_zz_255] <= _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port1 = RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0[_zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0];
  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port2 = RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0[_zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port_1) begin
      RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1[_zz_255] <= _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port1 = RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1[_zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0];
  assign _zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port2 = RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1[_zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_port) begin
      RobPlugin_logic_storage_BRANCH_HISTORY_banks_0[_zz_262] <= FrontendPlugin_allocated_BRANCH_HISTORY_0;
    end
  end

  assign _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_port1 = RobPlugin_logic_storage_BRANCH_HISTORY_banks_0[_zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_1_port) begin
      RobPlugin_logic_storage_BRANCH_HISTORY_banks_1[_zz_262] <= FrontendPlugin_allocated_BRANCH_HISTORY_1;
    end
  end

  assign _zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_1_port1 = RobPlugin_logic_storage_BRANCH_HISTORY_banks_1[_zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port_1) begin
      RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0[_zz_267] <= _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port1 = RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0[_zz_DecoderPredictionPlugin_logic_ras_healPush];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1_port_1) begin
      RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1[_zz_267] <= _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1_port1 = RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1[_zz_DecoderPredictionPlugin_logic_ras_healPush];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port_2) begin
      RobPlugin_logic_storage_LQ_ALLOC_banks_0[_zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port] <= _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port_1;
    end
  end

  assign _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port1 = RobPlugin_logic_storage_LQ_ALLOC_banks_0[_zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port_2) begin
      RobPlugin_logic_storage_SQ_ALLOC_banks_0[_zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port] <= _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port_1;
    end
  end

  assign _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port1 = RobPlugin_logic_storage_SQ_ALLOC_banks_0[_zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port) begin
      RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0[_zz_276] <= FrontendPlugin_allocated_Frontend_MICRO_OP_0;
    end
  end

  assign _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port1 = RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP];
  assign _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port2 = RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1_port) begin
      RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1[_zz_276] <= FrontendPlugin_allocated_Frontend_MICRO_OP_1;
    end
  end

  assign _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1_port1 = RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1[_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP];
  assign _zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1_port2 = RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port_1) begin
      RobPlugin_logic_storage_PHYS_RS_0_banks_0[_zz_283] <= _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_0_port1 = RobPlugin_logic_storage_PHYS_RS_0_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RS_0_banks_1_port_1) begin
      RobPlugin_logic_storage_PHYS_RS_0_banks_1[_zz_283] <= _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_PHYS_RS_0_banks_1_port1 = RobPlugin_logic_storage_PHYS_RS_0_banks_1[_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port_1) begin
      RobPlugin_logic_storage_READ_RS_0_banks_0[_zz_288] <= _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port1 = RobPlugin_logic_storage_READ_RS_0_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0];
  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port2 = RobPlugin_logic_storage_READ_RS_0_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port_1) begin
      RobPlugin_logic_storage_READ_RS_0_banks_1[_zz_288] <= _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port1 = RobPlugin_logic_storage_READ_RS_0_banks_1[_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0];
  assign _zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port2 = RobPlugin_logic_storage_READ_RS_0_banks_1[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port_1) begin
      RobPlugin_logic_storage_PHYS_RS_1_banks_0[_zz_295] <= _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_0_port1 = RobPlugin_logic_storage_PHYS_RS_1_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_PHYS_RS_1_banks_1_port_1) begin
      RobPlugin_logic_storage_PHYS_RS_1_banks_1[_zz_295] <= _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_PHYS_RS_1_banks_1_port1 = RobPlugin_logic_storage_PHYS_RS_1_banks_1[_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port_1) begin
      RobPlugin_logic_storage_READ_RS_1_banks_0[_zz_300] <= _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port1 = RobPlugin_logic_storage_READ_RS_1_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1];
  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port2 = RobPlugin_logic_storage_READ_RS_1_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port_1) begin
      RobPlugin_logic_storage_READ_RS_1_banks_1[_zz_300] <= _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port1 = RobPlugin_logic_storage_READ_RS_1_banks_1[_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1];
  assign _zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port2 = RobPlugin_logic_storage_READ_RS_1_banks_1[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port_1) begin
      RobPlugin_logic_storage_BRANCH_ID_banks_0[_zz_307] <= _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_BRANCH_ID_banks_0_port1 = RobPlugin_logic_storage_BRANCH_ID_banks_0[_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_BRANCH_ID_banks_1_port_1) begin
      RobPlugin_logic_storage_BRANCH_ID_banks_1[_zz_307] <= _zz_RobPlugin_logic_storage_BRANCH_ID_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_BRANCH_ID_banks_1_port1 = RobPlugin_logic_storage_BRANCH_ID_banks_1[_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_LSU_ID_banks_0_port_1) begin
      RobPlugin_logic_storage_LSU_ID_banks_0[_zz_312] <= _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_LSU_ID_banks_0_port1 = RobPlugin_logic_storage_LSU_ID_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_LSU_ID_banks_1_port_1) begin
      RobPlugin_logic_storage_LSU_ID_banks_1[_zz_312] <= _zz_RobPlugin_logic_storage_LSU_ID_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_LSU_ID_banks_1_port1 = RobPlugin_logic_storage_LSU_ID_banks_1[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port_1) begin
      RobPlugin_logic_storage_ROB_MSB_banks_0[_zz_317] <= _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port1 = RobPlugin_logic_storage_ROB_MSB_banks_0[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB];
  always @(posedge clk) begin
    if(_zz_RobPlugin_logic_storage_ROB_MSB_banks_1_port_1) begin
      RobPlugin_logic_storage_ROB_MSB_banks_1[_zz_317] <= _zz_RobPlugin_logic_storage_ROB_MSB_banks_1_port;
    end
  end

  assign _zz_RobPlugin_logic_storage_ROB_MSB_banks_1_port1 = RobPlugin_logic_storage_ROB_MSB_banks_1[_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB];
  TranslatorWithRollback integer_RfTranslationPlugin_logic_impl (
    .io_rollback                  (integer_RfTranslationPlugin_logic_impl_io_rollback                      ), //i
    .io_writes_0_valid            (integer_RfTranslationPlugin_logic_impl_io_writes_0_valid                ), //i
    .io_writes_0_payload_address  (FrontendPlugin_allocated_ARCH_RD_0[4:0]                                 ), //i
    .io_writes_0_payload_data     (FrontendPlugin_allocated_PHYS_RD_0[5:0]                                 ), //i
    .io_writes_1_valid            (integer_RfTranslationPlugin_logic_impl_io_writes_1_valid                ), //i
    .io_writes_1_payload_address  (FrontendPlugin_allocated_ARCH_RD_1[4:0]                                 ), //i
    .io_writes_1_payload_data     (FrontendPlugin_allocated_PHYS_RD_1[5:0]                                 ), //i
    .io_commits_0_valid           (integer_RfTranslationPlugin_logic_impl_io_commits_0_valid               ), //i
    .io_commits_0_payload_address (integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_address[4:0]), //i
    .io_commits_0_payload_data    (integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_data[5:0]   ), //i
    .io_commits_1_valid           (integer_RfTranslationPlugin_logic_impl_io_commits_1_valid               ), //i
    .io_commits_1_payload_address (integer_RfTranslationPlugin_logic_onCommit_archRd_1[4:0]                ), //i
    .io_commits_1_payload_data    (integer_RfTranslationPlugin_logic_onCommit_physRd_1[5:0]                ), //i
    .io_reads_0_cmd_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_0_cmd_valid             ), //i
    .io_reads_0_cmd_payload       (FrontendPlugin_allocated_ARCH_RD_0[4:0]                                 ), //i
    .io_reads_0_rsp_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_valid             ), //o
    .io_reads_0_rsp_payload       (integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_payload[5:0]      ), //o
    .io_reads_1_cmd_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_1_cmd_valid             ), //i
    .io_reads_1_cmd_payload       (FrontendPlugin_allocated_ARCH_RS_0_0[4:0]                               ), //i
    .io_reads_1_rsp_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_valid             ), //o
    .io_reads_1_rsp_payload       (integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_payload[5:0]      ), //o
    .io_reads_2_cmd_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_2_cmd_valid             ), //i
    .io_reads_2_cmd_payload       (FrontendPlugin_allocated_ARCH_RS_1_0[4:0]                               ), //i
    .io_reads_2_rsp_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_valid             ), //o
    .io_reads_2_rsp_payload       (integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_payload[5:0]      ), //o
    .io_reads_3_cmd_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_3_cmd_valid             ), //i
    .io_reads_3_cmd_payload       (FrontendPlugin_allocated_ARCH_RD_1[4:0]                                 ), //i
    .io_reads_3_rsp_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_3_rsp_valid             ), //o
    .io_reads_3_rsp_payload       (integer_RfTranslationPlugin_logic_impl_io_reads_3_rsp_payload[5:0]      ), //o
    .io_reads_4_cmd_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_4_cmd_valid             ), //i
    .io_reads_4_cmd_payload       (FrontendPlugin_allocated_ARCH_RS_0_1[4:0]                               ), //i
    .io_reads_4_rsp_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_4_rsp_valid             ), //o
    .io_reads_4_rsp_payload       (integer_RfTranslationPlugin_logic_impl_io_reads_4_rsp_payload[5:0]      ), //o
    .io_reads_5_cmd_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_5_cmd_valid             ), //i
    .io_reads_5_cmd_payload       (FrontendPlugin_allocated_ARCH_RS_1_1[4:0]                               ), //i
    .io_reads_5_rsp_valid         (integer_RfTranslationPlugin_logic_impl_io_reads_5_rsp_valid             ), //o
    .io_reads_5_rsp_payload       (integer_RfTranslationPlugin_logic_impl_io_reads_5_rsp_payload[5:0]      ), //o
    .clk                          (clk                                                                     ), //i
    .reset                        (reset                                                                   )  //i
  );
  AllocatorMultiPortMem integer_RfAllocationPlugin_logic_allocator (
    .io_push_0_valid   (integer_RfAllocationPlugin_logic_allocator_io_push_0_valid       ), //i
    .io_push_0_payload (integer_RfAllocationPlugin_logic_allocator_io_push_0_payload[5:0]), //i
    .io_push_1_valid   (integer_RfAllocationPlugin_logic_allocator_io_push_1_valid       ), //i
    .io_push_1_payload (integer_RfAllocationPlugin_logic_allocator_io_push_1_payload[5:0]), //i
    .io_pop_mask       (integer_RfAllocationPlugin_logic_allocator_io_pop_mask[1:0]      ), //i
    .io_pop_ready      (integer_RfAllocationPlugin_logic_allocator_io_pop_ready          ), //o
    .io_pop_fire       (FrontendPlugin_allocated_isFireing                               ), //i
    .io_pop_values_0   (integer_RfAllocationPlugin_logic_allocator_io_pop_values_0[5:0]  ), //o
    .io_pop_values_1   (integer_RfAllocationPlugin_logic_allocator_io_pop_values_1[5:0]  ), //o
    .clk               (clk                                                              ), //i
    .reset             (reset                                                            )  //i
  );
  DataCache DataCachePlugin_logic_cache (
    .io_lock_valid                             (DataCachePlugin_setup_lockPort_valid                                       ), //i
    .io_lock_address                           (DataCachePlugin_setup_lockPort_address[31:0]                               ), //i
    .io_load_cmd_valid                         (DataCachePlugin_logic_load_hit                                             ), //i
    .io_load_cmd_ready                         (DataCachePlugin_logic_cache_io_load_cmd_ready                              ), //o
    .io_load_cmd_payload_virtual               (DataCachePlugin_logic_cache_io_load_cmd_payload_virtual[31:0]              ), //i
    .io_load_cmd_payload_size                  (DataCachePlugin_logic_cache_io_load_cmd_payload_size[1:0]                  ), //i
    .io_load_cmd_payload_redoOnDataHazard      (DataCachePlugin_logic_cache_io_load_cmd_payload_redoOnDataHazard           ), //i
    .io_load_cmd_payload_unlocked              (DataCachePlugin_logic_cache_io_load_cmd_payload_unlocked                   ), //i
    .io_load_cmd_payload_unique                (DataCachePlugin_logic_cache_io_load_cmd_payload_unique                     ), //i
    .io_load_translated_physical               (DataCachePlugin_logic_cache_io_load_translated_physical[31:0]              ), //i
    .io_load_translated_abord                  (DataCachePlugin_logic_cache_io_load_translated_abord                       ), //i
    .io_load_cancels                           (DataCachePlugin_logic_cache_io_load_cancels[2:0]                           ), //i
    .io_load_rsp_valid                         (DataCachePlugin_logic_cache_io_load_rsp_valid                              ), //o
    .io_load_rsp_payload_data                  (DataCachePlugin_logic_cache_io_load_rsp_payload_data[31:0]                 ), //o
    .io_load_rsp_payload_fault                 (DataCachePlugin_logic_cache_io_load_rsp_payload_fault                      ), //o
    .io_load_rsp_payload_redo                  (DataCachePlugin_logic_cache_io_load_rsp_payload_redo                       ), //o
    .io_load_rsp_payload_refillSlot            (DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlot[1:0]            ), //o
    .io_load_rsp_payload_refillSlotAny         (DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlotAny              ), //o
    .io_store_cmd_valid                        (Lsu2Plugin_setup_cacheStore_cmd_valid                                      ), //i
    .io_store_cmd_ready                        (DataCachePlugin_logic_cache_io_store_cmd_ready                             ), //o
    .io_store_cmd_payload_address              (Lsu2Plugin_setup_cacheStore_cmd_payload_address[31:0]                      ), //i
    .io_store_cmd_payload_data                 (Lsu2Plugin_setup_cacheStore_cmd_payload_data[31:0]                         ), //i
    .io_store_cmd_payload_mask                 (Lsu2Plugin_setup_cacheStore_cmd_payload_mask[3:0]                          ), //i
    .io_store_cmd_payload_generation           (Lsu2Plugin_setup_cacheStore_cmd_payload_generation                         ), //i
    .io_store_cmd_payload_io                   (Lsu2Plugin_setup_cacheStore_cmd_payload_io                                 ), //i
    .io_store_cmd_payload_flush                (Lsu2Plugin_setup_cacheStore_cmd_payload_flush                              ), //i
    .io_store_cmd_payload_flushFree            (Lsu2Plugin_setup_cacheStore_cmd_payload_flushFree                          ), //i
    .io_store_cmd_payload_prefetch             (Lsu2Plugin_setup_cacheStore_cmd_payload_prefetch                           ), //i
    .io_store_rsp_valid                        (DataCachePlugin_logic_cache_io_store_rsp_valid                             ), //o
    .io_store_rsp_payload_fault                (DataCachePlugin_logic_cache_io_store_rsp_payload_fault                     ), //o
    .io_store_rsp_payload_redo                 (DataCachePlugin_logic_cache_io_store_rsp_payload_redo                      ), //o
    .io_store_rsp_payload_refillSlot           (DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlot[1:0]           ), //o
    .io_store_rsp_payload_refillSlotAny        (DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlotAny             ), //o
    .io_store_rsp_payload_generationKo         (DataCachePlugin_logic_cache_io_store_rsp_payload_generationKo              ), //o
    .io_store_rsp_payload_flush                (DataCachePlugin_logic_cache_io_store_rsp_payload_flush                     ), //o
    .io_store_rsp_payload_prefetch             (DataCachePlugin_logic_cache_io_store_rsp_payload_prefetch                  ), //o
    .io_store_rsp_payload_address              (DataCachePlugin_logic_cache_io_store_rsp_payload_address[31:0]             ), //o
    .io_store_rsp_payload_io                   (DataCachePlugin_logic_cache_io_store_rsp_payload_io                        ), //o
    .io_mem_read_cmd_valid                     (DataCachePlugin_logic_cache_io_mem_read_cmd_valid                          ), //o
    .io_mem_read_cmd_ready                     (DataCachePlugin_mem_read_cmd_ready                                         ), //i
    .io_mem_read_cmd_payload_id                (DataCachePlugin_logic_cache_io_mem_read_cmd_payload_id                     ), //o
    .io_mem_read_cmd_payload_address           (DataCachePlugin_logic_cache_io_mem_read_cmd_payload_address[31:0]          ), //o
    .io_mem_read_rsp_valid                     (DataCachePlugin_mem_read_rsp_valid                                         ), //i
    .io_mem_read_rsp_ready                     (DataCachePlugin_logic_cache_io_mem_read_rsp_ready                          ), //o
    .io_mem_read_rsp_payload_id                (DataCachePlugin_mem_read_rsp_payload_id                                    ), //i
    .io_mem_read_rsp_payload_data              (DataCachePlugin_mem_read_rsp_payload_data[63:0]                            ), //i
    .io_mem_read_rsp_payload_error             (DataCachePlugin_mem_read_rsp_payload_error                                 ), //i
    .io_mem_write_cmd_valid                    (DataCachePlugin_logic_cache_io_mem_write_cmd_valid                         ), //o
    .io_mem_write_cmd_ready                    (DataCachePlugin_mem_write_cmd_ready                                        ), //i
    .io_mem_write_cmd_payload_last             (DataCachePlugin_logic_cache_io_mem_write_cmd_payload_last                  ), //o
    .io_mem_write_cmd_payload_fragment_address (DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_address[31:0]), //o
    .io_mem_write_cmd_payload_fragment_data    (DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_data[63:0]   ), //o
    .io_mem_write_cmd_payload_fragment_id      (DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_id           ), //o
    .io_mem_write_rsp_valid                    (DataCachePlugin_mem_write_rsp_valid                                        ), //i
    .io_mem_write_rsp_payload_error            (DataCachePlugin_mem_write_rsp_payload_error                                ), //i
    .io_mem_write_rsp_payload_id               (DataCachePlugin_mem_write_rsp_payload_id                                   ), //i
    .io_refillCompletions                      (DataCachePlugin_logic_cache_io_refillCompletions[1:0]                      ), //o
    .io_refillEvent                            (DataCachePlugin_logic_cache_io_refillEvent                                 ), //o
    .io_writebackEvent                         (DataCachePlugin_logic_cache_io_writebackEvent                              ), //o
    .io_writebackBusy                          (DataCachePlugin_logic_cache_io_writebackBusy                               ), //o
    .io_tagEvent                               (DataCachePlugin_logic_cache_io_tagEvent                                    ), //o
    .clk                                       (clk                                                                        ), //i
    .reset                                     (reset                                                                      )  //i
  );
  StreamFifoLowLatency CommitPlugin_logic_free_lineEventStream_fifo (
    .io_push_valid         (CommitPlugin_logic_free_lineEventStream_valid                         ), //i
    .io_push_ready         (CommitPlugin_logic_free_lineEventStream_fifo_io_push_ready            ), //o
    .io_push_payload_robId (CommitPlugin_logic_free_lineEventStream_payload_robId[5:0]            ), //i
    .io_push_payload_mask  (CommitPlugin_logic_free_lineEventStream_payload_mask[1:0]             ), //i
    .io_pop_valid          (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_valid             ), //o
    .io_pop_ready          (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_ready             ), //i
    .io_pop_payload_robId  (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_robId[5:0]), //o
    .io_pop_payload_mask   (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_mask[1:0] ), //o
    .io_flush              (CommitPlugin_logic_free_lineEventStream_fifo_io_flush                 ), //i
    .io_occupancy          (CommitPlugin_logic_free_lineEventStream_fifo_io_occupancy[5:0]        ), //o
    .io_availability       (CommitPlugin_logic_free_lineEventStream_fifo_io_availability[5:0]     ), //o
    .clk                   (clk                                                                   ), //i
    .reset                 (reset                                                                 )  //i
  );
  DivRadix4 EU0_DivPlugin_logic_div (
    .io_flush              (EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed                          ), //i
    .io_cmd_valid          (EU0_DivPlugin_logic_div_io_cmd_valid                                        ), //i
    .io_cmd_ready          (EU0_DivPlugin_logic_div_io_cmd_ready                                        ), //o
    .io_cmd_payload_a      (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED[31:0]), //i
    .io_cmd_payload_b      (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED[31:0]), //i
    .io_rsp_valid          (EU0_DivPlugin_logic_div_io_rsp_valid                                        ), //o
    .io_rsp_ready          (EU0_ExecutionUnitBase_pipeline_execute_1_ready                              ), //i
    .io_rsp_payload_result (EU0_DivPlugin_logic_div_io_rsp_payload_result[34:0]                         ), //o
    .io_rsp_payload_remain (EU0_DivPlugin_logic_div_io_rsp_payload_remain[32:0]                         ), //o
    .clk                   (clk                                                                         ), //i
    .reset                 (reset                                                                       )  //i
  );
  PrefetchPredictor Lsu2Plugin_logic_prefetch_predictor (
    .io_learn_valid            (Lsu2Plugin_logic_prefetch_predictor_io_learn_valid                 ), //i
    .io_learn_payload_physical (Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_address[31:0]     ), //i
    .io_learn_payload_allocate (Lsu2Plugin_logic_prefetch_predictor_io_learn_payload_allocate      ), //i
    .io_prediction_cmd_valid   (Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_valid        ), //o
    .io_prediction_cmd_ready   (Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready        ), //i
    .io_prediction_cmd_payload (Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_payload[31:0]), //o
    .io_prediction_rsp_valid   (Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_valid        ), //i
    .io_prediction_rsp_payload (Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_payload      )  //i
  );
  IssueQueue DispatchPlugin_logic_queue (
    .io_clear                                   (CommitPlugin_logic_commit_reschedulePort_valid                       ), //i
    .io_events                                  (DispatchPlugin_logic_wake_optReduce_reduced[31:0]                    ), //i
    .io_push_valid                              (FrontendPlugin_dispatch_isFireing                                    ), //i
    .io_push_ready                              (DispatchPlugin_logic_queue_io_push_ready                             ), //o
    .io_push_payload_slots_0_event              (DispatchPlugin_logic_queue_io_push_payload_slots_0_event[31:0]       ), //i
    .io_push_payload_slots_0_sel                (DispatchPlugin_logic_queue_io_push_payload_slots_0_sel[1:0]          ), //i
    .io_push_payload_slots_0_context_staticWake (DispatchPlugin_logic_queue_io_push_payload_slots_0_context_staticWake), //i
    .io_push_payload_slots_0_context_physRd     (FrontendPlugin_dispatch_PHYS_RD_0[5:0]                               ), //i
    .io_push_payload_slots_0_context_robId      (DispatchPlugin_logic_queue_io_push_payload_slots_0_context_robId[5:0]), //i
    .io_push_payload_slots_0_context_euCtx_0    (FrontendPlugin_dispatch_PHYS_RS_0_0[5:0]                             ), //i
    .io_push_payload_slots_0_context_euCtx_1    (FrontendPlugin_dispatch_PHYS_RS_1_0[5:0]                             ), //i
    .io_push_payload_slots_1_event              (DispatchPlugin_logic_queue_io_push_payload_slots_1_event[31:0]       ), //i
    .io_push_payload_slots_1_sel                (DispatchPlugin_logic_queue_io_push_payload_slots_1_sel[1:0]          ), //i
    .io_push_payload_slots_1_context_staticWake (DispatchPlugin_logic_queue_io_push_payload_slots_1_context_staticWake), //i
    .io_push_payload_slots_1_context_physRd     (FrontendPlugin_dispatch_PHYS_RD_1[5:0]                               ), //i
    .io_push_payload_slots_1_context_robId      (DispatchPlugin_logic_queue_io_push_payload_slots_1_context_robId[5:0]), //i
    .io_push_payload_slots_1_context_euCtx_0    (FrontendPlugin_dispatch_PHYS_RS_0_1[5:0]                             ), //i
    .io_push_payload_slots_1_context_euCtx_1    (FrontendPlugin_dispatch_PHYS_RS_1_1[5:0]                             ), //i
    .io_schedules_0_valid                       (DispatchPlugin_logic_queue_io_schedules_0_valid                      ), //o
    .io_schedules_0_ready                       (DispatchPlugin_logic_pop_0_stagesList_0_ready                        ), //i
    .io_schedules_0_payload_event               (DispatchPlugin_logic_queue_io_schedules_0_payload_event[15:0]        ), //o
    .io_schedules_1_valid                       (DispatchPlugin_logic_queue_io_schedules_1_valid                      ), //o
    .io_schedules_1_ready                       (DispatchPlugin_logic_pop_1_stagesList_0_ready                        ), //i
    .io_schedules_1_payload_event               (DispatchPlugin_logic_queue_io_schedules_1_payload_event[15:0]        ), //o
    .io_schedules_2_valid                       (DispatchPlugin_logic_queue_io_schedules_2_valid                      ), //o
    .io_schedules_2_ready                       (DispatchPlugin_logic_pop_2_stagesList_0_ready                        ), //i
    .io_schedules_2_payload_event               (DispatchPlugin_logic_queue_io_schedules_2_payload_event[31:0]        ), //o
    .io_contexts_0_staticWake                   (DispatchPlugin_logic_queue_io_contexts_0_staticWake                  ), //o
    .io_contexts_0_physRd                       (DispatchPlugin_logic_queue_io_contexts_0_physRd[5:0]                 ), //o
    .io_contexts_0_robId                        (DispatchPlugin_logic_queue_io_contexts_0_robId[5:0]                  ), //o
    .io_contexts_0_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_0_euCtx_0[5:0]                ), //o
    .io_contexts_0_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_0_euCtx_1[5:0]                ), //o
    .io_contexts_1_staticWake                   (DispatchPlugin_logic_queue_io_contexts_1_staticWake                  ), //o
    .io_contexts_1_physRd                       (DispatchPlugin_logic_queue_io_contexts_1_physRd[5:0]                 ), //o
    .io_contexts_1_robId                        (DispatchPlugin_logic_queue_io_contexts_1_robId[5:0]                  ), //o
    .io_contexts_1_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_1_euCtx_0[5:0]                ), //o
    .io_contexts_1_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_1_euCtx_1[5:0]                ), //o
    .io_contexts_2_staticWake                   (DispatchPlugin_logic_queue_io_contexts_2_staticWake                  ), //o
    .io_contexts_2_physRd                       (DispatchPlugin_logic_queue_io_contexts_2_physRd[5:0]                 ), //o
    .io_contexts_2_robId                        (DispatchPlugin_logic_queue_io_contexts_2_robId[5:0]                  ), //o
    .io_contexts_2_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_2_euCtx_0[5:0]                ), //o
    .io_contexts_2_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_2_euCtx_1[5:0]                ), //o
    .io_contexts_3_staticWake                   (DispatchPlugin_logic_queue_io_contexts_3_staticWake                  ), //o
    .io_contexts_3_physRd                       (DispatchPlugin_logic_queue_io_contexts_3_physRd[5:0]                 ), //o
    .io_contexts_3_robId                        (DispatchPlugin_logic_queue_io_contexts_3_robId[5:0]                  ), //o
    .io_contexts_3_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_3_euCtx_0[5:0]                ), //o
    .io_contexts_3_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_3_euCtx_1[5:0]                ), //o
    .io_contexts_4_staticWake                   (DispatchPlugin_logic_queue_io_contexts_4_staticWake                  ), //o
    .io_contexts_4_physRd                       (DispatchPlugin_logic_queue_io_contexts_4_physRd[5:0]                 ), //o
    .io_contexts_4_robId                        (DispatchPlugin_logic_queue_io_contexts_4_robId[5:0]                  ), //o
    .io_contexts_4_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_4_euCtx_0[5:0]                ), //o
    .io_contexts_4_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_4_euCtx_1[5:0]                ), //o
    .io_contexts_5_staticWake                   (DispatchPlugin_logic_queue_io_contexts_5_staticWake                  ), //o
    .io_contexts_5_physRd                       (DispatchPlugin_logic_queue_io_contexts_5_physRd[5:0]                 ), //o
    .io_contexts_5_robId                        (DispatchPlugin_logic_queue_io_contexts_5_robId[5:0]                  ), //o
    .io_contexts_5_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_5_euCtx_0[5:0]                ), //o
    .io_contexts_5_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_5_euCtx_1[5:0]                ), //o
    .io_contexts_6_staticWake                   (DispatchPlugin_logic_queue_io_contexts_6_staticWake                  ), //o
    .io_contexts_6_physRd                       (DispatchPlugin_logic_queue_io_contexts_6_physRd[5:0]                 ), //o
    .io_contexts_6_robId                        (DispatchPlugin_logic_queue_io_contexts_6_robId[5:0]                  ), //o
    .io_contexts_6_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_6_euCtx_0[5:0]                ), //o
    .io_contexts_6_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_6_euCtx_1[5:0]                ), //o
    .io_contexts_7_staticWake                   (DispatchPlugin_logic_queue_io_contexts_7_staticWake                  ), //o
    .io_contexts_7_physRd                       (DispatchPlugin_logic_queue_io_contexts_7_physRd[5:0]                 ), //o
    .io_contexts_7_robId                        (DispatchPlugin_logic_queue_io_contexts_7_robId[5:0]                  ), //o
    .io_contexts_7_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_7_euCtx_0[5:0]                ), //o
    .io_contexts_7_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_7_euCtx_1[5:0]                ), //o
    .io_contexts_8_staticWake                   (DispatchPlugin_logic_queue_io_contexts_8_staticWake                  ), //o
    .io_contexts_8_physRd                       (DispatchPlugin_logic_queue_io_contexts_8_physRd[5:0]                 ), //o
    .io_contexts_8_robId                        (DispatchPlugin_logic_queue_io_contexts_8_robId[5:0]                  ), //o
    .io_contexts_8_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_8_euCtx_0[5:0]                ), //o
    .io_contexts_8_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_8_euCtx_1[5:0]                ), //o
    .io_contexts_9_staticWake                   (DispatchPlugin_logic_queue_io_contexts_9_staticWake                  ), //o
    .io_contexts_9_physRd                       (DispatchPlugin_logic_queue_io_contexts_9_physRd[5:0]                 ), //o
    .io_contexts_9_robId                        (DispatchPlugin_logic_queue_io_contexts_9_robId[5:0]                  ), //o
    .io_contexts_9_euCtx_0                      (DispatchPlugin_logic_queue_io_contexts_9_euCtx_0[5:0]                ), //o
    .io_contexts_9_euCtx_1                      (DispatchPlugin_logic_queue_io_contexts_9_euCtx_1[5:0]                ), //o
    .io_contexts_10_staticWake                  (DispatchPlugin_logic_queue_io_contexts_10_staticWake                 ), //o
    .io_contexts_10_physRd                      (DispatchPlugin_logic_queue_io_contexts_10_physRd[5:0]                ), //o
    .io_contexts_10_robId                       (DispatchPlugin_logic_queue_io_contexts_10_robId[5:0]                 ), //o
    .io_contexts_10_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_10_euCtx_0[5:0]               ), //o
    .io_contexts_10_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_10_euCtx_1[5:0]               ), //o
    .io_contexts_11_staticWake                  (DispatchPlugin_logic_queue_io_contexts_11_staticWake                 ), //o
    .io_contexts_11_physRd                      (DispatchPlugin_logic_queue_io_contexts_11_physRd[5:0]                ), //o
    .io_contexts_11_robId                       (DispatchPlugin_logic_queue_io_contexts_11_robId[5:0]                 ), //o
    .io_contexts_11_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_11_euCtx_0[5:0]               ), //o
    .io_contexts_11_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_11_euCtx_1[5:0]               ), //o
    .io_contexts_12_staticWake                  (DispatchPlugin_logic_queue_io_contexts_12_staticWake                 ), //o
    .io_contexts_12_physRd                      (DispatchPlugin_logic_queue_io_contexts_12_physRd[5:0]                ), //o
    .io_contexts_12_robId                       (DispatchPlugin_logic_queue_io_contexts_12_robId[5:0]                 ), //o
    .io_contexts_12_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_12_euCtx_0[5:0]               ), //o
    .io_contexts_12_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_12_euCtx_1[5:0]               ), //o
    .io_contexts_13_staticWake                  (DispatchPlugin_logic_queue_io_contexts_13_staticWake                 ), //o
    .io_contexts_13_physRd                      (DispatchPlugin_logic_queue_io_contexts_13_physRd[5:0]                ), //o
    .io_contexts_13_robId                       (DispatchPlugin_logic_queue_io_contexts_13_robId[5:0]                 ), //o
    .io_contexts_13_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_13_euCtx_0[5:0]               ), //o
    .io_contexts_13_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_13_euCtx_1[5:0]               ), //o
    .io_contexts_14_staticWake                  (DispatchPlugin_logic_queue_io_contexts_14_staticWake                 ), //o
    .io_contexts_14_physRd                      (DispatchPlugin_logic_queue_io_contexts_14_physRd[5:0]                ), //o
    .io_contexts_14_robId                       (DispatchPlugin_logic_queue_io_contexts_14_robId[5:0]                 ), //o
    .io_contexts_14_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_14_euCtx_0[5:0]               ), //o
    .io_contexts_14_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_14_euCtx_1[5:0]               ), //o
    .io_contexts_15_staticWake                  (DispatchPlugin_logic_queue_io_contexts_15_staticWake                 ), //o
    .io_contexts_15_physRd                      (DispatchPlugin_logic_queue_io_contexts_15_physRd[5:0]                ), //o
    .io_contexts_15_robId                       (DispatchPlugin_logic_queue_io_contexts_15_robId[5:0]                 ), //o
    .io_contexts_15_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_15_euCtx_0[5:0]               ), //o
    .io_contexts_15_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_15_euCtx_1[5:0]               ), //o
    .io_contexts_16_staticWake                  (DispatchPlugin_logic_queue_io_contexts_16_staticWake                 ), //o
    .io_contexts_16_physRd                      (DispatchPlugin_logic_queue_io_contexts_16_physRd[5:0]                ), //o
    .io_contexts_16_robId                       (DispatchPlugin_logic_queue_io_contexts_16_robId[5:0]                 ), //o
    .io_contexts_16_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_16_euCtx_0[5:0]               ), //o
    .io_contexts_16_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_16_euCtx_1[5:0]               ), //o
    .io_contexts_17_staticWake                  (DispatchPlugin_logic_queue_io_contexts_17_staticWake                 ), //o
    .io_contexts_17_physRd                      (DispatchPlugin_logic_queue_io_contexts_17_physRd[5:0]                ), //o
    .io_contexts_17_robId                       (DispatchPlugin_logic_queue_io_contexts_17_robId[5:0]                 ), //o
    .io_contexts_17_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_17_euCtx_0[5:0]               ), //o
    .io_contexts_17_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_17_euCtx_1[5:0]               ), //o
    .io_contexts_18_staticWake                  (DispatchPlugin_logic_queue_io_contexts_18_staticWake                 ), //o
    .io_contexts_18_physRd                      (DispatchPlugin_logic_queue_io_contexts_18_physRd[5:0]                ), //o
    .io_contexts_18_robId                       (DispatchPlugin_logic_queue_io_contexts_18_robId[5:0]                 ), //o
    .io_contexts_18_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_18_euCtx_0[5:0]               ), //o
    .io_contexts_18_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_18_euCtx_1[5:0]               ), //o
    .io_contexts_19_staticWake                  (DispatchPlugin_logic_queue_io_contexts_19_staticWake                 ), //o
    .io_contexts_19_physRd                      (DispatchPlugin_logic_queue_io_contexts_19_physRd[5:0]                ), //o
    .io_contexts_19_robId                       (DispatchPlugin_logic_queue_io_contexts_19_robId[5:0]                 ), //o
    .io_contexts_19_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_19_euCtx_0[5:0]               ), //o
    .io_contexts_19_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_19_euCtx_1[5:0]               ), //o
    .io_contexts_20_staticWake                  (DispatchPlugin_logic_queue_io_contexts_20_staticWake                 ), //o
    .io_contexts_20_physRd                      (DispatchPlugin_logic_queue_io_contexts_20_physRd[5:0]                ), //o
    .io_contexts_20_robId                       (DispatchPlugin_logic_queue_io_contexts_20_robId[5:0]                 ), //o
    .io_contexts_20_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_20_euCtx_0[5:0]               ), //o
    .io_contexts_20_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_20_euCtx_1[5:0]               ), //o
    .io_contexts_21_staticWake                  (DispatchPlugin_logic_queue_io_contexts_21_staticWake                 ), //o
    .io_contexts_21_physRd                      (DispatchPlugin_logic_queue_io_contexts_21_physRd[5:0]                ), //o
    .io_contexts_21_robId                       (DispatchPlugin_logic_queue_io_contexts_21_robId[5:0]                 ), //o
    .io_contexts_21_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_21_euCtx_0[5:0]               ), //o
    .io_contexts_21_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_21_euCtx_1[5:0]               ), //o
    .io_contexts_22_staticWake                  (DispatchPlugin_logic_queue_io_contexts_22_staticWake                 ), //o
    .io_contexts_22_physRd                      (DispatchPlugin_logic_queue_io_contexts_22_physRd[5:0]                ), //o
    .io_contexts_22_robId                       (DispatchPlugin_logic_queue_io_contexts_22_robId[5:0]                 ), //o
    .io_contexts_22_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_22_euCtx_0[5:0]               ), //o
    .io_contexts_22_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_22_euCtx_1[5:0]               ), //o
    .io_contexts_23_staticWake                  (DispatchPlugin_logic_queue_io_contexts_23_staticWake                 ), //o
    .io_contexts_23_physRd                      (DispatchPlugin_logic_queue_io_contexts_23_physRd[5:0]                ), //o
    .io_contexts_23_robId                       (DispatchPlugin_logic_queue_io_contexts_23_robId[5:0]                 ), //o
    .io_contexts_23_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_23_euCtx_0[5:0]               ), //o
    .io_contexts_23_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_23_euCtx_1[5:0]               ), //o
    .io_contexts_24_staticWake                  (DispatchPlugin_logic_queue_io_contexts_24_staticWake                 ), //o
    .io_contexts_24_physRd                      (DispatchPlugin_logic_queue_io_contexts_24_physRd[5:0]                ), //o
    .io_contexts_24_robId                       (DispatchPlugin_logic_queue_io_contexts_24_robId[5:0]                 ), //o
    .io_contexts_24_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_24_euCtx_0[5:0]               ), //o
    .io_contexts_24_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_24_euCtx_1[5:0]               ), //o
    .io_contexts_25_staticWake                  (DispatchPlugin_logic_queue_io_contexts_25_staticWake                 ), //o
    .io_contexts_25_physRd                      (DispatchPlugin_logic_queue_io_contexts_25_physRd[5:0]                ), //o
    .io_contexts_25_robId                       (DispatchPlugin_logic_queue_io_contexts_25_robId[5:0]                 ), //o
    .io_contexts_25_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_25_euCtx_0[5:0]               ), //o
    .io_contexts_25_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_25_euCtx_1[5:0]               ), //o
    .io_contexts_26_staticWake                  (DispatchPlugin_logic_queue_io_contexts_26_staticWake                 ), //o
    .io_contexts_26_physRd                      (DispatchPlugin_logic_queue_io_contexts_26_physRd[5:0]                ), //o
    .io_contexts_26_robId                       (DispatchPlugin_logic_queue_io_contexts_26_robId[5:0]                 ), //o
    .io_contexts_26_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_26_euCtx_0[5:0]               ), //o
    .io_contexts_26_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_26_euCtx_1[5:0]               ), //o
    .io_contexts_27_staticWake                  (DispatchPlugin_logic_queue_io_contexts_27_staticWake                 ), //o
    .io_contexts_27_physRd                      (DispatchPlugin_logic_queue_io_contexts_27_physRd[5:0]                ), //o
    .io_contexts_27_robId                       (DispatchPlugin_logic_queue_io_contexts_27_robId[5:0]                 ), //o
    .io_contexts_27_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_27_euCtx_0[5:0]               ), //o
    .io_contexts_27_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_27_euCtx_1[5:0]               ), //o
    .io_contexts_28_staticWake                  (DispatchPlugin_logic_queue_io_contexts_28_staticWake                 ), //o
    .io_contexts_28_physRd                      (DispatchPlugin_logic_queue_io_contexts_28_physRd[5:0]                ), //o
    .io_contexts_28_robId                       (DispatchPlugin_logic_queue_io_contexts_28_robId[5:0]                 ), //o
    .io_contexts_28_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_28_euCtx_0[5:0]               ), //o
    .io_contexts_28_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_28_euCtx_1[5:0]               ), //o
    .io_contexts_29_staticWake                  (DispatchPlugin_logic_queue_io_contexts_29_staticWake                 ), //o
    .io_contexts_29_physRd                      (DispatchPlugin_logic_queue_io_contexts_29_physRd[5:0]                ), //o
    .io_contexts_29_robId                       (DispatchPlugin_logic_queue_io_contexts_29_robId[5:0]                 ), //o
    .io_contexts_29_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_29_euCtx_0[5:0]               ), //o
    .io_contexts_29_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_29_euCtx_1[5:0]               ), //o
    .io_contexts_30_staticWake                  (DispatchPlugin_logic_queue_io_contexts_30_staticWake                 ), //o
    .io_contexts_30_physRd                      (DispatchPlugin_logic_queue_io_contexts_30_physRd[5:0]                ), //o
    .io_contexts_30_robId                       (DispatchPlugin_logic_queue_io_contexts_30_robId[5:0]                 ), //o
    .io_contexts_30_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_30_euCtx_0[5:0]               ), //o
    .io_contexts_30_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_30_euCtx_1[5:0]               ), //o
    .io_contexts_31_staticWake                  (DispatchPlugin_logic_queue_io_contexts_31_staticWake                 ), //o
    .io_contexts_31_physRd                      (DispatchPlugin_logic_queue_io_contexts_31_physRd[5:0]                ), //o
    .io_contexts_31_robId                       (DispatchPlugin_logic_queue_io_contexts_31_robId[5:0]                 ), //o
    .io_contexts_31_euCtx_0                     (DispatchPlugin_logic_queue_io_contexts_31_euCtx_0[5:0]               ), //o
    .io_contexts_31_euCtx_1                     (DispatchPlugin_logic_queue_io_contexts_31_euCtx_1[5:0]               ), //o
    .io_usage                                   (DispatchPlugin_logic_queue_io_usage[31:0]                            ), //o
    .clk                                        (clk                                                                  ), //i
    .reset                                      (reset                                                                )  //i
  );
  RegFileAsync integer_RegFilePlugin_logic_regfile_fpga (
    .io_writes_0_valid   (integer_RegFilePlugin_logic_writeMerges_0_bus_valid             ), //i
    .io_writes_0_address (integer_RegFilePlugin_logic_writeMerges_0_bus_address[5:0]      ), //i
    .io_writes_0_data    (integer_RegFilePlugin_logic_writeMerges_0_bus_data[31:0]        ), //i
    .io_writes_0_robId   (integer_RegFilePlugin_logic_writeMerges_0_bus_robId[5:0]        ), //i
    .io_writes_1_valid   (integer_RegFilePlugin_logic_writeMerges_1_bus_valid             ), //i
    .io_writes_1_address (integer_RegFilePlugin_logic_writeMerges_1_bus_address[5:0]      ), //i
    .io_writes_1_data    (integer_RegFilePlugin_logic_writeMerges_1_bus_data[31:0]        ), //i
    .io_writes_1_robId   (integer_RegFilePlugin_logic_writeMerges_1_bus_robId[5:0]        ), //i
    .io_writes_2_valid   (integer_RegFilePlugin_logic_writeMerges_2_bus_valid             ), //i
    .io_writes_2_address (integer_RegFilePlugin_logic_writeMerges_2_bus_address[5:0]      ), //i
    .io_writes_2_data    (integer_RegFilePlugin_logic_writeMerges_2_bus_data[31:0]        ), //i
    .io_writes_2_robId   (integer_RegFilePlugin_logic_writeMerges_2_bus_robId[5:0]        ), //i
    .io_writes_3_valid   (integer_RegFilePlugin_logic_writeMerges_3_bus_valid             ), //i
    .io_writes_3_address (integer_RegFilePlugin_logic_writeMerges_3_bus_address[5:0]      ), //i
    .io_writes_3_data    (integer_RegFilePlugin_logic_writeMerges_3_bus_data[31:0]        ), //i
    .io_writes_3_robId   (integer_RegFilePlugin_logic_writeMerges_3_bus_robId[5:0]        ), //i
    .io_reads_0_valid    (ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid       ), //i
    .io_reads_0_address  (ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address[5:0]), //i
    .io_reads_0_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data[31:0]  ), //o
    .io_reads_1_valid    (ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid       ), //i
    .io_reads_1_address  (ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address[5:0]), //i
    .io_reads_1_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data[31:0]  ), //o
    .io_reads_2_valid    (ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid       ), //i
    .io_reads_2_address  (ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address[5:0]), //i
    .io_reads_2_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_2_data[31:0]  ), //o
    .io_reads_3_valid    (ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid       ), //i
    .io_reads_3_address  (ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address[5:0]), //i
    .io_reads_3_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_3_data[31:0]  ), //o
    .io_reads_4_valid    (EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid        ), //i
    .io_reads_4_address  (EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address[5:0] ), //i
    .io_reads_4_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_4_data[31:0]  ), //o
    .io_reads_5_valid    (EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid        ), //i
    .io_reads_5_address  (EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address[5:0] ), //i
    .io_reads_5_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_5_data[31:0]  ), //o
    .clk                 (clk                                                             ), //i
    .reset               (reset                                                           )  //i
  );
  DependencyStorage RfDependencyPlugin_logic_forRf_integer_impl (
    .io_writes_0_valid             (RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_valid                 ), //i
    .io_writes_0_payload_physical  (FrontendPlugin_dispatch_PHYS_RD_0[5:0]                                        ), //i
    .io_writes_0_payload_robId     (RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_payload_robId[5:0]    ), //i
    .io_writes_1_valid             (RfDependencyPlugin_logic_forRf_integer_impl_io_writes_1_valid                 ), //i
    .io_writes_1_payload_physical  (FrontendPlugin_dispatch_PHYS_RD_1[5:0]                                        ), //i
    .io_writes_1_payload_robId     (RfDependencyPlugin_logic_forRf_integer_impl_io_writes_1_payload_robId[5:0]    ), //i
    .io_commits_0_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_valid                ), //i
    .io_commits_0_payload_physical (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_payload_physical[5:0]), //i
    .io_commits_1_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_1_valid                ), //i
    .io_commits_1_payload_physical (DispatchPlugin_logic_pop_1_wake_L0_bypassed_payload_physical[5:0]             ), //i
    .io_commits_2_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_2_valid                ), //i
    .io_commits_2_payload_physical (Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_payload_physical[5:0]        ), //i
    .io_commits_3_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_3_valid                ), //i
    .io_commits_3_payload_physical (Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_payload_physical[5:0]                  ), //i
    .io_commits_4_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_4_valid                ), //i
    .io_commits_4_payload_physical (Lsu2Plugin_logic_special_wakeRf_payload_physical[5:0]                         ), //i
    .io_commits_5_valid            (RfDependencyPlugin_logic_forRf_integer_impl_io_commits_5_valid                ), //i
    .io_commits_5_payload_physical (EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_payload_physical[5:0]        ), //i
    .io_reads_0_cmd_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_cmd_valid              ), //i
    .io_reads_0_cmd_payload        (FrontendPlugin_dispatch_PHYS_RS_0_0[5:0]                                      ), //i
    .io_reads_0_rsp_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_valid              ), //o
    .io_reads_0_rsp_payload_enable (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_enable     ), //o
    .io_reads_0_rsp_payload_rob    (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_rob[5:0]   ), //o
    .io_reads_1_cmd_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_cmd_valid              ), //i
    .io_reads_1_cmd_payload        (FrontendPlugin_dispatch_PHYS_RS_1_0[5:0]                                      ), //i
    .io_reads_1_rsp_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_valid              ), //o
    .io_reads_1_rsp_payload_enable (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_enable     ), //o
    .io_reads_1_rsp_payload_rob    (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_rob[5:0]   ), //o
    .io_reads_2_cmd_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_cmd_valid              ), //i
    .io_reads_2_cmd_payload        (FrontendPlugin_dispatch_PHYS_RS_0_1[5:0]                                      ), //i
    .io_reads_2_rsp_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_rsp_valid              ), //o
    .io_reads_2_rsp_payload_enable (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_rsp_payload_enable     ), //o
    .io_reads_2_rsp_payload_rob    (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_rsp_payload_rob[5:0]   ), //o
    .io_reads_3_cmd_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_cmd_valid              ), //i
    .io_reads_3_cmd_payload        (FrontendPlugin_dispatch_PHYS_RS_1_1[5:0]                                      ), //i
    .io_reads_3_rsp_valid          (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_rsp_valid              ), //o
    .io_reads_3_rsp_payload_enable (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_rsp_payload_enable     ), //o
    .io_reads_3_rsp_payload_rob    (RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_rsp_payload_rob[5:0]   ), //o
    .clk                           (clk                                                                           ), //i
    .reset                         (reset                                                                         )  //i
  );
  RamAsyncMwMux BranchContextPlugin_logic_mem_earlyBranch (
    .io_writes_0_valid           (_zz_io_writes_0_valid_7                                                 ), //i
    .io_writes_0_payload_address (FrontendPlugin_allocated_BRANCH_ID_0[3:0]                               ), //i
    .io_writes_0_payload_data    (BranchContextPlugin_logic_mem_earlyBranch_io_writes_0_payload_data[32:0]), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid_9                                                 ), //i
    .io_writes_1_payload_address (FrontendPlugin_allocated_BRANCH_ID_1[3:0]                               ), //i
    .io_writes_1_payload_data    (BranchContextPlugin_logic_mem_earlyBranch_io_writes_1_payload_data[32:0]), //i
    .io_read_0_cmd_valid         (BranchContextPlugin_logic_mem_earlyBranch_io_read_0_cmd_valid           ), //i
    .io_read_0_cmd_payload       (ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID[3:0]                ), //i
    .io_read_0_rsp               (BranchContextPlugin_logic_mem_earlyBranch_io_read_0_rsp[32:0]           ), //o
    .io_read_1_cmd_valid         (BranchContextPlugin_logic_mem_earlyBranch_io_read_1_cmd_valid           ), //i
    .io_read_1_cmd_payload       (ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID[3:0]                ), //i
    .io_read_1_rsp               (BranchContextPlugin_logic_mem_earlyBranch_io_read_1_rsp[32:0]           ), //o
    .clk                         (clk                                                                     ), //i
    .reset                       (reset                                                                   )  //i
  );
  RamAsyncMwMux_1 BranchContextPlugin_logic_mem_finalBranch (
    .io_writes_0_valid           (_zz_io_writes_0_valid_1                                                 ), //i
    .io_writes_0_payload_address (ALU0_BranchPlugin_logic_branch_finalBranch_payload_address[3:0]         ), //i
    .io_writes_0_payload_data    (BranchContextPlugin_logic_mem_finalBranch_io_writes_0_payload_data[64:0]), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid_1                                                 ), //i
    .io_writes_1_payload_address (ALU1_BranchPlugin_logic_branch_finalBranch_payload_address[3:0]         ), //i
    .io_writes_1_payload_data    (BranchContextPlugin_logic_mem_finalBranch_io_writes_1_payload_data[64:0]), //i
    .io_read_0_cmd_valid         (BranchContextPlugin_logic_mem_finalBranch_io_read_0_cmd_valid           ), //i
    .io_read_0_cmd_payload       (BranchContextPlugin_free_learn_bid[3:0]                                 ), //i
    .io_read_0_rsp               (BranchContextPlugin_logic_mem_finalBranch_io_read_0_rsp[64:0]           ), //o
    .clk                         (clk                                                                     ), //i
    .reset                       (reset                                                                   )  //i
  );
  RamAsyncMwXor Lsu2Plugin_logic_lq_mem_sqAlloc (
    .io_writes_0_valid           (_zz_io_writes_0_valid_6                                      ), //i
    .io_writes_0_payload_address (FrontendPlugin_dispatch_LQ_ID_0[3:0]                         ), //i
    .io_writes_0_payload_data    (Lsu2Plugin_logic_lq_mem_sqAlloc_io_writes_0_payload_data[4:0]), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid_8                                      ), //i
    .io_writes_1_payload_address (FrontendPlugin_dispatch_LQ_ID_1[3:0]                         ), //i
    .io_writes_1_payload_data    (Lsu2Plugin_logic_lq_mem_sqAlloc_io_writes_1_payload_data[4:0]), //i
    .io_read_0_cmd_valid         (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_0_cmd_valid          ), //i
    .io_read_0_cmd_payload       (Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID[3:0]               ), //i
    .io_read_0_rsp               (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_0_rsp[4:0]           ), //o
    .io_read_1_cmd_valid         (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_1_cmd_valid          ), //i
    .io_read_1_cmd_payload       (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_1_cmd_payload[3:0]   ), //i
    .io_read_1_rsp               (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_1_rsp[4:0]           ), //o
    .io_read_2_cmd_valid         (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_2_cmd_valid          ), //i
    .io_read_2_cmd_payload       (Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID[3:0]               ), //i
    .io_read_2_rsp               (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_2_rsp[4:0]           ), //o
    .io_read_3_cmd_valid         (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_3_cmd_valid          ), //i
    .io_read_3_cmd_payload       (Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ID[3:0]     ), //i
    .io_read_3_rsp               (Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_3_rsp[4:0]           ), //o
    .clk                         (clk                                                          ), //i
    .reset                       (reset                                                        )  //i
  );
  RamAsyncMwXor_1 Lsu2Plugin_logic_lq_mem_doSpecial (
    .io_writes_0_valid           (_zz_io_writes_0_valid_5                                   ), //i
    .io_writes_0_payload_address (FrontendPlugin_dispatch_LQ_ID_0[3:0]                      ), //i
    .io_writes_0_payload_data    (Lsu2Plugin_logic_lq_mem_doSpecial_io_writes_0_payload_data), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid_7                                   ), //i
    .io_writes_1_payload_address (FrontendPlugin_dispatch_LQ_ID_1[3:0]                      ), //i
    .io_writes_1_payload_data    (Lsu2Plugin_logic_lq_mem_doSpecial_io_writes_1_payload_data), //i
    .io_writes_2_valid           (_zz_io_writes_2_valid_1                                   ), //i
    .io_writes_2_payload_address (Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID[3:0]            ), //i
    .io_writes_2_payload_data    (Lsu2Plugin_logic_lq_mem_doSpecial_io_writes_2_payload_data), //i
    .io_read_0_cmd_valid         (Lsu2Plugin_logic_lq_mem_doSpecial_io_read_0_cmd_valid     ), //i
    .io_read_0_cmd_payload       (Lsu2Plugin_logic_lq_ptr_freeReal[3:0]                     ), //i
    .io_read_0_rsp               (Lsu2Plugin_logic_lq_mem_doSpecial_io_read_0_rsp           ), //o
    .clk                         (clk                                                       ), //i
    .reset                       (reset                                                     )  //i
  );
  RamAsyncMwXor_9 Lsu2Plugin_logic_lq_mem_needTranslation (
    .io_writes_0_valid           (Lsu2Plugin_logic_aguPush_0_pushLq                                       ), //i
    .io_writes_0_payload_address (Lsu2Plugin_logic_lq_mem_needTranslation_io_writes_0_payload_address[3:0]), //i
    .io_writes_0_payload_data    (Lsu2Plugin_logic_lq_mem_needTranslation_io_writes_0_payload_data        ), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid_3                                                 ), //i
    .io_writes_1_payload_address (Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID[3:0]                          ), //i
    .io_writes_1_payload_data    (Lsu2Plugin_logic_lq_mem_needTranslation_io_writes_1_payload_data        ), //i
    .io_read_0_cmd_valid         (Lsu2Plugin_logic_lq_mem_needTranslation_io_read_0_cmd_valid             ), //i
    .io_read_0_cmd_payload       (Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID[3:0]                          ), //i
    .io_read_0_rsp               (Lsu2Plugin_logic_lq_mem_needTranslation_io_read_0_rsp                   ), //o
    .clk                         (clk                                                                     ), //i
    .reset                       (reset                                                                   )  //i
  );
  RamAsyncMwXor_10 Lsu2Plugin_logic_sq_mem_needTranslation (
    .io_writes_0_valid           (Lsu2Plugin_logic_aguPush_0_pushSq                                       ), //i
    .io_writes_0_payload_address (Lsu2Plugin_logic_sq_mem_needTranslation_io_writes_0_payload_address[3:0]), //i
    .io_writes_0_payload_data    (Lsu2Plugin_logic_sq_mem_needTranslation_io_writes_0_payload_data        ), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid_2                                                 ), //i
    .io_writes_1_payload_address (Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID[3:0]                          ), //i
    .io_writes_1_payload_data    (Lsu2Plugin_logic_sq_mem_needTranslation_io_writes_1_payload_data        ), //i
    .io_read_0_cmd_valid         (Lsu2Plugin_logic_sq_mem_needTranslation_io_read_0_cmd_valid             ), //i
    .io_read_0_cmd_payload       (Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID[3:0]                          ), //i
    .io_read_0_rsp               (Lsu2Plugin_logic_sq_mem_needTranslation_io_read_0_rsp                   ), //o
    .io_read_1_cmd_valid         (Lsu2Plugin_logic_sq_mem_needTranslation_io_read_1_cmd_valid             ), //i
    .io_read_1_cmd_payload       (Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID[3:0]                 ), //i
    .io_read_1_rsp               (Lsu2Plugin_logic_sq_mem_needTranslation_io_read_1_rsp                   ), //o
    .clk                         (clk                                                                     ), //i
    .reset                       (reset                                                                   )  //i
  );
  RamAsyncMwXor_1 Lsu2Plugin_logic_sq_mem_feededOnce (
    .io_writes_0_valid           (_zz_io_writes_0_valid_2                                       ), //i
    .io_writes_0_payload_address (FrontendPlugin_dispatch_SQ_ID_0[3:0]                          ), //i
    .io_writes_0_payload_data    (Lsu2Plugin_logic_sq_mem_feededOnce_io_writes_0_payload_data   ), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid_4                                       ), //i
    .io_writes_1_payload_address (FrontendPlugin_dispatch_SQ_ID_1[3:0]                          ), //i
    .io_writes_1_payload_data    (Lsu2Plugin_logic_sq_mem_feededOnce_io_writes_1_payload_data   ), //i
    .io_writes_2_valid           (_zz_io_writes_2_valid_2                                       ), //i
    .io_writes_2_payload_address (Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID[3:0]                ), //i
    .io_writes_2_payload_data    (Lsu2Plugin_logic_sq_mem_feededOnce_io_writes_2_payload_data   ), //i
    .io_read_0_cmd_valid         (Lsu2Plugin_logic_sq_mem_feededOnce_io_read_0_cmd_valid        ), //i
    .io_read_0_cmd_payload       (Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SQID[3:0]), //i
    .io_read_0_rsp               (Lsu2Plugin_logic_sq_mem_feededOnce_io_read_0_rsp              ), //o
    .clk                         (clk                                                           ), //i
    .reset                       (reset                                                         )  //i
  );
  RamAsyncMwXor_1 Lsu2Plugin_logic_sq_mem_doSpecial (
    .io_writes_0_valid           (_zz_io_writes_0_valid_4                                   ), //i
    .io_writes_0_payload_address (FrontendPlugin_dispatch_SQ_ID_0[3:0]                      ), //i
    .io_writes_0_payload_data    (Lsu2Plugin_logic_sq_mem_doSpecial_io_writes_0_payload_data), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid_6                                   ), //i
    .io_writes_1_payload_address (FrontendPlugin_dispatch_SQ_ID_1[3:0]                      ), //i
    .io_writes_1_payload_data    (Lsu2Plugin_logic_sq_mem_doSpecial_io_writes_1_payload_data), //i
    .io_writes_2_valid           (_zz_io_writes_2_valid                                     ), //i
    .io_writes_2_payload_address (Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID[3:0]            ), //i
    .io_writes_2_payload_data    (Lsu2Plugin_logic_sq_mem_doSpecial_io_writes_2_payload_data), //i
    .io_read_0_cmd_valid         (Lsu2Plugin_logic_sq_mem_doSpecial_io_read_0_cmd_valid     ), //i
    .io_read_0_cmd_payload       (Lsu2Plugin_logic_sq_ptr_commitReal[3:0]                   ), //i
    .io_read_0_rsp               (Lsu2Plugin_logic_sq_mem_doSpecial_io_read_0_rsp           ), //o
    .clk                         (clk                                                       ), //i
    .reset                       (reset                                                     )  //i
  );
  RamAsyncMwXor_6 Lsu2Plugin_logic_sq_mem_lqAlloc (
    .io_writes_0_valid           (_zz_io_writes_0_valid_3                                      ), //i
    .io_writes_0_payload_address (FrontendPlugin_dispatch_SQ_ID_0[3:0]                         ), //i
    .io_writes_0_payload_data    (Lsu2Plugin_logic_sq_mem_lqAlloc_io_writes_0_payload_data[4:0]), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid_5                                      ), //i
    .io_writes_1_payload_address (FrontendPlugin_dispatch_SQ_ID_1[3:0]                         ), //i
    .io_writes_1_payload_data    (Lsu2Plugin_logic_sq_mem_lqAlloc_io_writes_1_payload_data[4:0]), //i
    .io_read_0_cmd_valid         (Lsu2Plugin_logic_sq_mem_lqAlloc_io_read_0_cmd_valid          ), //i
    .io_read_0_cmd_payload       (Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID[3:0]               ), //i
    .io_read_0_rsp               (Lsu2Plugin_logic_sq_mem_lqAlloc_io_read_0_rsp[4:0]           ), //o
    .clk                         (clk                                                          ), //i
    .reset                       (reset                                                        )  //i
  );
  RamAsyncMwMux_2 BranchContextPlugin_free_dispatchMem_mem (
    .io_writes_0_valid           (_zz_io_writes_0_valid                                                  ), //i
    .io_writes_0_payload_address (BranchContextPlugin_free_dispatchMem_writes_0_port_payload_address[3:0]), //i
    .io_writes_0_payload_data    (BranchContextPlugin_free_dispatchMem_writes_0_port_payload_data[28:0]  ), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid                                                  ), //i
    .io_writes_1_payload_address (BranchContextPlugin_free_dispatchMem_writes_1_port_payload_address[3:0]), //i
    .io_writes_1_payload_data    (BranchContextPlugin_free_dispatchMem_writes_1_port_payload_data[28:0]  ), //i
    .io_read_0_cmd_valid         (BranchContextPlugin_free_dispatchMem_mem_io_read_0_cmd_valid           ), //i
    .io_read_0_cmd_payload       (BranchContextPlugin_free_learn_bid[3:0]                                ), //i
    .io_read_0_rsp               (BranchContextPlugin_free_dispatchMem_mem_io_read_0_rsp[28:0]           ), //o
    .clk                         (clk                                                                    ), //i
    .reset                       (reset                                                                  )  //i
  );
  RamAsyncMwXor_7 RobPlugin_logic_storage_BRANCH_TAKEN_banks_0 (
    .io_writes_0_valid           (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_0_valid         ), //i
    .io_writes_0_payload_address (ALU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID[5:0]                  ), //i
    .io_writes_0_payload_data    (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_0_payload_data  ), //i
    .io_writes_1_valid           (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_1_valid         ), //i
    .io_writes_1_payload_address (ALU1_ExecutionUnitBase_pipeline_execute_1_ROB_ID[5:0]                  ), //i
    .io_writes_1_payload_data    (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_1_payload_data  ), //i
    .io_read_0_cmd_valid         (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_0_cmd_valid       ), //i
    .io_read_0_cmd_payload       (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_0_cmd_payload[5:0]), //i
    .io_read_0_rsp               (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_0_rsp             ), //o
    .io_read_1_cmd_valid         (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_1_cmd_valid       ), //i
    .io_read_1_cmd_payload       (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_1_cmd_payload[5:0]), //i
    .io_read_1_rsp               (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_1_rsp             ), //o
    .io_read_2_cmd_valid         (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_2_cmd_valid       ), //i
    .io_read_2_cmd_payload       (CommitPlugin_logic_reschedule_reschedulePort_payload_robId[5:0]        ), //i
    .io_read_2_rsp               (RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_2_rsp             ), //o
    .clk                         (clk                                                                    ), //i
    .reset                       (reset                                                                  )  //i
  );
  always @(*) begin
    case(_zz_FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT_1)
      1'b0 : _zz_FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT = 2'b11;
      default : _zz_FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT = 2'b10;
    endcase
  end

  always @(*) begin
    case(AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_SLICE)
      1'b0 : _zz_AlignerPlugin_setup_s2m_MASK_BACK = 2'b01;
      default : _zz_AlignerPlugin_setup_s2m_MASK_BACK = 2'b11;
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_extractors_0_pcWord_1)
      1'b0 : _zz_AlignerPlugin_logic_extractors_0_pcWord = AlignerPlugin_logic_buffer_pc;
      default : _zz_AlignerPlugin_logic_extractors_0_pcWord = AlignerPlugin_setup_s2m_Fetch_FETCH_PC;
    endcase
  end

  always @(*) begin
    case(_zz_AlignerPlugin_logic_extractors_1_pcWord_1)
      1'b0 : _zz_AlignerPlugin_logic_extractors_1_pcWord = AlignerPlugin_logic_buffer_pc;
      default : _zz_AlignerPlugin_logic_extractors_1_pcWord = AlignerPlugin_setup_s2m_Fetch_FETCH_PC;
    endcase
  end

  always @(*) begin
    case(FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_slice)
      1'b0 : _zz_BtbPlugin_logic_applyIt_prediction = FetchPlugin_stages_1_GSHARE_COUNTER_0[1];
      default : _zz_BtbPlugin_logic_applyIt_prediction = FetchPlugin_stages_1_GSHARE_COUNTER_1[1];
    endcase
  end

  always @(*) begin
    case(_zz_CommitDebugFilterPlugin_logic_commits_3)
      2'b00 : _zz_CommitDebugFilterPlugin_logic_commits_2 = 2'b00;
      2'b01 : _zz_CommitDebugFilterPlugin_logic_commits_2 = 2'b01;
      2'b10 : _zz_CommitDebugFilterPlugin_logic_commits_2 = 2'b01;
      default : _zz_CommitDebugFilterPlugin_logic_commits_2 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_3)
      1'b0 : _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_2 = _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_1[31 : 0];
      default : _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_2 = _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_1[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_commitCount_1)
      2'b00 : _zz_PerformanceCounterPlugin_logic_commitCount = 2'b00;
      2'b01 : _zz_PerformanceCounterPlugin_logic_commitCount = 2'b01;
      2'b10 : _zz_PerformanceCounterPlugin_logic_commitCount = 2'b01;
      default : _zz_PerformanceCounterPlugin_logic_commitCount = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_0_1)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_0 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_0 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_1_1)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_2_1)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_2 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_2 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_3_1)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_3 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_3 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_BranchContextPlugin_logic_onCommit_commitedNext_2)
      2'b00 : _zz_BranchContextPlugin_logic_onCommit_commitedNext_1 = 2'b00;
      2'b01 : _zz_BranchContextPlugin_logic_onCommit_commitedNext_1 = 2'b01;
      2'b10 : _zz_BranchContextPlugin_logic_onCommit_commitedNext_1 = 2'b01;
      default : _zz_BranchContextPlugin_logic_onCommit_commitedNext_1 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_3)
      1'b0 : _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_2 = _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_1[23 : 0];
      default : _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_2 = _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_1[47 : 24];
    endcase
  end

  always @(*) begin
    case(_zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_3)
      1'b0 : _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_2 = _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_1[0 : 0];
      default : _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_2 = _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_1[1 : 1];
    endcase
  end

  always @(*) begin
    case(_zz_DecoderPredictionPlugin_logic_ras_healPush_3)
      1'b0 : _zz_DecoderPredictionPlugin_logic_ras_healPush_2 = _zz_DecoderPredictionPlugin_logic_ras_healPush_1[3 : 0];
      default : _zz_DecoderPredictionPlugin_logic_ras_healPush_2 = _zz_DecoderPredictionPlugin_logic_ras_healPush_1[7 : 4];
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount_1)
      2'b00 : _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount = 2'b00;
      2'b01 : _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount = 2'b01;
      2'b10 : _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount = 2'b01;
      default : _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_allocation_loads_requestsCount_1)
      2'b00 : _zz_Lsu2Plugin_logic_allocation_loads_requestsCount = 2'b00;
      2'b01 : _zz_Lsu2Plugin_logic_allocation_loads_requestsCount = 2'b01;
      2'b10 : _zz_Lsu2Plugin_logic_allocation_loads_requestsCount = 2'b01;
      default : _zz_Lsu2Plugin_logic_allocation_loads_requestsCount = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_allocation_stores_requestsCount_1)
      2'b00 : _zz_Lsu2Plugin_logic_allocation_stores_requestsCount = 2'b00;
      2'b01 : _zz_Lsu2Plugin_logic_allocation_stores_requestsCount = 2'b01;
      2'b10 : _zz_Lsu2Plugin_logic_allocation_stores_requestsCount = 2'b01;
      default : _zz_Lsu2Plugin_logic_allocation_stores_requestsCount = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_1)
      2'b00 : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_0;
      2'b01 : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_1;
      2'b10 : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_2;
      default : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3;
    endcase
  end

  always @(*) begin
    case(_zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_3)
      1'b0 : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_2 = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_1;
      default : _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_2 = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3;
    endcase
  end

  always @(*) begin
    case(Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID)
      4'b0000 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_0_niceHazard;
      4'b0001 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_1_niceHazard;
      4'b0010 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_2_niceHazard;
      4'b0011 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_3_niceHazard;
      4'b0100 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_4_niceHazard;
      4'b0101 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_5_niceHazard;
      4'b0110 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_6_niceHazard;
      4'b0111 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_7_niceHazard;
      4'b1000 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_8_niceHazard;
      4'b1001 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_9_niceHazard;
      4'b1010 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_10_niceHazard;
      4'b1011 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_11_niceHazard;
      4'b1100 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_12_niceHazard;
      4'b1101 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_13_niceHazard;
      4'b1110 : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_14_niceHazard;
      default : _zz__zz_when_Lsu2Plugin_l1348 = Lsu2Plugin_logic_lq_regs_15_niceHazard;
    endcase
  end

  always @(*) begin
    case(CsrRamPlugin_logic_writeLogic_sel)
      2'b00 : begin
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_address = EU0_CsrAccessPlugin_logic_ramWritePort_address;
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_data = EU0_CsrAccessPlugin_logic_ramWritePort_data;
      end
      2'b01 : begin
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_address = PerformanceCounterPlugin_setup_writePort_address;
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_data = PerformanceCounterPlugin_setup_writePort_data;
      end
      2'b10 : begin
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_address = PrivilegedPlugin_setup_ramWrite_address;
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_data = PrivilegedPlugin_setup_ramWrite_data;
      end
      default : begin
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_address = CsrRamPlugin_setup_initPort_address;
        _zz_CsrRamPlugin_logic_writeLogic_port_payload_data = CsrRamPlugin_setup_initPort_data;
      end
    endcase
  end

  always @(*) begin
    case(CsrRamPlugin_logic_readLogic_sel)
      2'b00 : _zz_CsrRamPlugin_logic_readLogic_port_address = EU0_CsrAccessPlugin_logic_ramReadPort_address;
      2'b01 : _zz_CsrRamPlugin_logic_readLogic_port_address = PerformanceCounterPlugin_setup_readPort_address;
      default : _zz_CsrRamPlugin_logic_readLogic_port_address = PrivilegedPlugin_setup_ramRead_address;
    endcase
  end

  always @(*) begin
    case(_zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17_1)
      1'b0 : _zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 = PerformanceCounterPlugin_logic_fsm_resultCsr[31 : 0];
      default : _zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 = PerformanceCounterPlugin_logic_fsm_resultCsr[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_3)
      1'b0 : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1[31 : 0];
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_3)
      1'b0 : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1[0 : 0];
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1[1 : 1];
    endcase
  end

  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_3)
      1'b0 : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1[0 : 0];
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1[1 : 1];
    endcase
  end

  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_3)
      1'b0 : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1[0 : 0];
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1[1 : 1];
    endcase
  end

  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_3)
      1'b0 : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_1[31 : 0];
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_1[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_3)
      1'b0 : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_1[4 : 0];
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_1[9 : 5];
    endcase
  end

  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_3)
      1'b0 : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_1[0 : 0];
      default : _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_1[1 : 1];
    endcase
  end

  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_3)
      2'b00 : _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2 = integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data;
      2'b01 : _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2 = integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data;
      default : _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2 = integer_RegFilePlugin_logic_writeMerges_2_bypass_port_data;
    endcase
  end

  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_3)
      2'b00 : _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2 = integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data;
      2'b01 : _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2 = integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data;
      default : _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2 = integer_RegFilePlugin_logic_writeMerges_2_bypass_port_data;
    endcase
  end

  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_3)
      2'b00 : _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2 = integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data;
      2'b01 : _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2 = integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data;
      default : _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2 = integer_RegFilePlugin_logic_writeMerges_2_bypass_port_data;
    endcase
  end

  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_3)
      2'b00 : _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2 = integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data;
      2'b01 : _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2 = integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data;
      default : _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2 = integer_RegFilePlugin_logic_writeMerges_2_bypass_port_data;
    endcase
  end

  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_3)
      2'b00 : _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2 = integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data;
      2'b01 : _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2 = integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data;
      default : _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2 = integer_RegFilePlugin_logic_writeMerges_2_bypass_port_data;
    endcase
  end

  always @(*) begin
    case(_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_3)
      2'b00 : _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2 = integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data;
      2'b01 : _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2 = integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data;
      default : _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2 = integer_RegFilePlugin_logic_writeMerges_2_bypass_port_data;
    endcase
  end

  always @(*) begin
    case(PerformanceCounterPlugin_logic_fsm_cmd_address)
      3'b000 : _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_11 = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded;
      3'b001 : _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_11 = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_1;
      3'b010 : _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_11 = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2;
      3'b011 : _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_11 = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3;
      3'b100 : _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_11 = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4;
      3'b101 : _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_11 = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5;
      default : _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_11 = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
      Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "TRAP_ALIGN ";
      Lsu2Plugin_CTRL_ENUM_MMU_REDO : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "MMU_REDO   ";
      Lsu2Plugin_CTRL_ENUM_TRAP_MMU : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "TRAP_MMU   ";
      Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "LOAD_HAZARD";
      Lsu2Plugin_CTRL_ENUM_LOAD_MISS : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "LOAD_MISS  ";
      Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "LOAD_FAILED";
      Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "TRAP_ACCESS";
      Lsu2Plugin_CTRL_ENUM_SUCCESS : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "SUCCESS    ";
      default : Lsu2Plugin_logic_sharedPip_stages_3_CTRL_string = "???????????";
    endcase
  end
  always @(*) begin
    case(Lsu2Plugin_logic_sharedPip_stages_2_CTRL)
      Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "TRAP_ALIGN ";
      Lsu2Plugin_CTRL_ENUM_MMU_REDO : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "MMU_REDO   ";
      Lsu2Plugin_CTRL_ENUM_TRAP_MMU : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "TRAP_MMU   ";
      Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "LOAD_HAZARD";
      Lsu2Plugin_CTRL_ENUM_LOAD_MISS : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "LOAD_MISS  ";
      Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "LOAD_FAILED";
      Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "TRAP_ACCESS";
      Lsu2Plugin_CTRL_ENUM_SUCCESS : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "SUCCESS    ";
      default : Lsu2Plugin_logic_sharedPip_stages_2_CTRL_string = "???????????";
    endcase
  end
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_BOOT : EnvCallPlugin_logic_flushes_stateReg_string = "BOOT           ";
      EnvCallPlugin_logic_flushes_enumDef_IDLE : EnvCallPlugin_logic_flushes_stateReg_string = "IDLE           ";
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : EnvCallPlugin_logic_flushes_stateReg_string = "RESCHEDULE     ";
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : EnvCallPlugin_logic_flushes_stateReg_string = "VMA_FETCH_FLUSH";
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : EnvCallPlugin_logic_flushes_stateReg_string = "VMA_FETCH_WAIT ";
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : EnvCallPlugin_logic_flushes_stateReg_string = "LSU_FLUSH      ";
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : EnvCallPlugin_logic_flushes_stateReg_string = "WAIT_LSU       ";
      default : EnvCallPlugin_logic_flushes_stateReg_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(EnvCallPlugin_logic_flushes_stateNext)
      EnvCallPlugin_logic_flushes_enumDef_BOOT : EnvCallPlugin_logic_flushes_stateNext_string = "BOOT           ";
      EnvCallPlugin_logic_flushes_enumDef_IDLE : EnvCallPlugin_logic_flushes_stateNext_string = "IDLE           ";
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : EnvCallPlugin_logic_flushes_stateNext_string = "RESCHEDULE     ";
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : EnvCallPlugin_logic_flushes_stateNext_string = "VMA_FETCH_FLUSH";
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : EnvCallPlugin_logic_flushes_stateNext_string = "VMA_FETCH_WAIT ";
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : EnvCallPlugin_logic_flushes_stateNext_string = "LSU_FLUSH      ";
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : EnvCallPlugin_logic_flushes_stateNext_string = "WAIT_LSU       ";
      default : EnvCallPlugin_logic_flushes_stateNext_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(Lsu2Plugin_logic_special_atomic_stateReg)
      Lsu2Plugin_logic_special_atomic_enumDef_BOOT : Lsu2Plugin_logic_special_atomic_stateReg_string = "BOOT      ";
      Lsu2Plugin_logic_special_atomic_enumDef_IDLE : Lsu2Plugin_logic_special_atomic_stateReg_string = "IDLE      ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD : Lsu2Plugin_logic_special_atomic_stateReg_string = "LOAD_CMD  ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP : Lsu2Plugin_logic_special_atomic_stateReg_string = "LOAD_RSP  ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY : Lsu2Plugin_logic_special_atomic_stateReg_string = "LOCK_DELAY";
      Lsu2Plugin_logic_special_atomic_enumDef_ALU : Lsu2Plugin_logic_special_atomic_stateReg_string = "ALU       ";
      Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION : Lsu2Plugin_logic_special_atomic_stateReg_string = "COMPLETION";
      Lsu2Plugin_logic_special_atomic_enumDef_SYNC : Lsu2Plugin_logic_special_atomic_stateReg_string = "SYNC      ";
      Lsu2Plugin_logic_special_atomic_enumDef_TRAP : Lsu2Plugin_logic_special_atomic_stateReg_string = "TRAP      ";
      default : Lsu2Plugin_logic_special_atomic_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(Lsu2Plugin_logic_special_atomic_stateNext)
      Lsu2Plugin_logic_special_atomic_enumDef_BOOT : Lsu2Plugin_logic_special_atomic_stateNext_string = "BOOT      ";
      Lsu2Plugin_logic_special_atomic_enumDef_IDLE : Lsu2Plugin_logic_special_atomic_stateNext_string = "IDLE      ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD : Lsu2Plugin_logic_special_atomic_stateNext_string = "LOAD_CMD  ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP : Lsu2Plugin_logic_special_atomic_stateNext_string = "LOAD_RSP  ";
      Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY : Lsu2Plugin_logic_special_atomic_stateNext_string = "LOCK_DELAY";
      Lsu2Plugin_logic_special_atomic_enumDef_ALU : Lsu2Plugin_logic_special_atomic_stateNext_string = "ALU       ";
      Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION : Lsu2Plugin_logic_special_atomic_stateNext_string = "COMPLETION";
      Lsu2Plugin_logic_special_atomic_enumDef_SYNC : Lsu2Plugin_logic_special_atomic_stateNext_string = "SYNC      ";
      Lsu2Plugin_logic_special_atomic_enumDef_TRAP : Lsu2Plugin_logic_special_atomic_stateNext_string = "TRAP      ";
      default : Lsu2Plugin_logic_special_atomic_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_BOOT : MmuPlugin_logic_refill_stateReg_string = "BOOT ";
      MmuPlugin_logic_refill_enumDef_IDLE : MmuPlugin_logic_refill_stateReg_string = "IDLE ";
      MmuPlugin_logic_refill_enumDef_INIT : MmuPlugin_logic_refill_stateReg_string = "INIT ";
      MmuPlugin_logic_refill_enumDef_CMD_0 : MmuPlugin_logic_refill_stateReg_string = "CMD_0";
      MmuPlugin_logic_refill_enumDef_CMD_1 : MmuPlugin_logic_refill_stateReg_string = "CMD_1";
      MmuPlugin_logic_refill_enumDef_RSP_0 : MmuPlugin_logic_refill_stateReg_string = "RSP_0";
      MmuPlugin_logic_refill_enumDef_RSP_1 : MmuPlugin_logic_refill_stateReg_string = "RSP_1";
      default : MmuPlugin_logic_refill_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateNext)
      MmuPlugin_logic_refill_enumDef_BOOT : MmuPlugin_logic_refill_stateNext_string = "BOOT ";
      MmuPlugin_logic_refill_enumDef_IDLE : MmuPlugin_logic_refill_stateNext_string = "IDLE ";
      MmuPlugin_logic_refill_enumDef_INIT : MmuPlugin_logic_refill_stateNext_string = "INIT ";
      MmuPlugin_logic_refill_enumDef_CMD_0 : MmuPlugin_logic_refill_stateNext_string = "CMD_0";
      MmuPlugin_logic_refill_enumDef_CMD_1 : MmuPlugin_logic_refill_stateNext_string = "CMD_1";
      MmuPlugin_logic_refill_enumDef_RSP_0 : MmuPlugin_logic_refill_stateNext_string = "RSP_0";
      MmuPlugin_logic_refill_enumDef_RSP_1 : MmuPlugin_logic_refill_stateNext_string = "RSP_1";
      default : MmuPlugin_logic_refill_stateNext_string = "?????";
    endcase
  end
  always @(*) begin
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "BOOT ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "IDLE ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "READ ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "WRITE";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "DONE ";
      default : EU0_CsrAccessPlugin_logic_fsm_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(EU0_CsrAccessPlugin_logic_fsm_stateNext)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "BOOT ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "IDLE ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "READ ";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "WRITE";
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "DONE ";
      default : EU0_CsrAccessPlugin_logic_fsm_stateNext_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "BITWISE ";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "AND_1";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1)
      BranchPlugin_BranchCtrlEnum_B : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "JALR";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2)
      BranchPlugin_BranchCtrlEnum_B : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "JALR";
      default : _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "BITWISE ";
      default : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2)
      IntAluPlugin_AluCtrlEnum_ADD_SUB : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "ADD_SUB ";
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "SLT_SLTU";
      IntAluPlugin_AluCtrlEnum_BITWISE : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "BITWISE ";
      default : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "AND_1";
      default : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_B : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "JALR";
      default : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1)
      BranchPlugin_BranchCtrlEnum_B : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "JALR";
      default : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2)
      BranchPlugin_BranchCtrlEnum_B : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "JALR";
      default : _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2_string = "????";
    endcase
  end
  always @(*) begin
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_BOOT : PerformanceCounterPlugin_logic_fsm_stateReg_string = "BOOT                ";
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : PerformanceCounterPlugin_logic_fsm_stateReg_string = "IDLE                ";
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : PerformanceCounterPlugin_logic_fsm_stateReg_string = "READ_LOW            ";
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : PerformanceCounterPlugin_logic_fsm_stateReg_string = "CALC                ";
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : PerformanceCounterPlugin_logic_fsm_stateReg_string = "WRITE_LOW           ";
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : PerformanceCounterPlugin_logic_fsm_stateReg_string = "READ_HIGH           ";
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : PerformanceCounterPlugin_logic_fsm_stateReg_string = "WRITE_HIGH          ";
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : PerformanceCounterPlugin_logic_fsm_stateReg_string = "CSR_WRITE           ";
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : PerformanceCounterPlugin_logic_fsm_stateReg_string = "CSR_WRITE_COMPLETION";
      default : PerformanceCounterPlugin_logic_fsm_stateReg_string = "????????????????????";
    endcase
  end
  always @(*) begin
    case(PerformanceCounterPlugin_logic_fsm_stateNext)
      PerformanceCounterPlugin_logic_fsm_enumDef_BOOT : PerformanceCounterPlugin_logic_fsm_stateNext_string = "BOOT                ";
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : PerformanceCounterPlugin_logic_fsm_stateNext_string = "IDLE                ";
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : PerformanceCounterPlugin_logic_fsm_stateNext_string = "READ_LOW            ";
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : PerformanceCounterPlugin_logic_fsm_stateNext_string = "CALC                ";
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : PerformanceCounterPlugin_logic_fsm_stateNext_string = "WRITE_LOW           ";
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : PerformanceCounterPlugin_logic_fsm_stateNext_string = "READ_HIGH           ";
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : PerformanceCounterPlugin_logic_fsm_stateNext_string = "WRITE_HIGH          ";
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : PerformanceCounterPlugin_logic_fsm_stateNext_string = "CSR_WRITE           ";
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : PerformanceCounterPlugin_logic_fsm_stateNext_string = "CSR_WRITE_COMPLETION";
      default : PerformanceCounterPlugin_logic_fsm_stateNext_string = "????????????????????";
    endcase
  end
  always @(*) begin
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_BOOT : PrivilegedPlugin_logic_fsm_stateReg_string = "BOOT      ";
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : PrivilegedPlugin_logic_fsm_stateReg_string = "IDLE      ";
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : PrivilegedPlugin_logic_fsm_stateReg_string = "SETUP     ";
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : PrivilegedPlugin_logic_fsm_stateReg_string = "EPC_WRITE ";
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : PrivilegedPlugin_logic_fsm_stateReg_string = "TVAL_WRITE";
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : PrivilegedPlugin_logic_fsm_stateReg_string = "EPC_READ  ";
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : PrivilegedPlugin_logic_fsm_stateReg_string = "TVEC_READ ";
      PrivilegedPlugin_logic_fsm_enumDef_XRET : PrivilegedPlugin_logic_fsm_stateReg_string = "XRET      ";
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : PrivilegedPlugin_logic_fsm_stateReg_string = "FLUSH_CALC";
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : PrivilegedPlugin_logic_fsm_stateReg_string = "FLUSH_JUMP";
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : PrivilegedPlugin_logic_fsm_stateReg_string = "TRAP      ";
      default : PrivilegedPlugin_logic_fsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(PrivilegedPlugin_logic_fsm_stateNext)
      PrivilegedPlugin_logic_fsm_enumDef_BOOT : PrivilegedPlugin_logic_fsm_stateNext_string = "BOOT      ";
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : PrivilegedPlugin_logic_fsm_stateNext_string = "IDLE      ";
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : PrivilegedPlugin_logic_fsm_stateNext_string = "SETUP     ";
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : PrivilegedPlugin_logic_fsm_stateNext_string = "EPC_WRITE ";
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : PrivilegedPlugin_logic_fsm_stateNext_string = "TVAL_WRITE";
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : PrivilegedPlugin_logic_fsm_stateNext_string = "EPC_READ  ";
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : PrivilegedPlugin_logic_fsm_stateNext_string = "TVEC_READ ";
      PrivilegedPlugin_logic_fsm_enumDef_XRET : PrivilegedPlugin_logic_fsm_stateNext_string = "XRET      ";
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : PrivilegedPlugin_logic_fsm_stateNext_string = "FLUSH_CALC";
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : PrivilegedPlugin_logic_fsm_stateNext_string = "FLUSH_JUMP";
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : PrivilegedPlugin_logic_fsm_stateNext_string = "TRAP      ";
      default : PrivilegedPlugin_logic_fsm_stateNext_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    if(EU0_ExecutionUnitBase_pipeline_completion_0_port_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(ALU1_ExecutionUnitBase_pipeline_completion_1_port_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_3 = 1'b0;
    if(ALU1_ExecutionUnitBase_pipeline_completion_0_port_valid) begin
      _zz_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_4 = 1'b0;
    if(ALU0_ExecutionUnitBase_pipeline_completion_1_port_valid) begin
      _zz_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_5 = 1'b0;
    if(ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid) begin
      _zz_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_6 = 1'b0;
    if(Lsu2Plugin_setup_specialCompletion_valid) begin
      _zz_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_7 = 1'b0;
    if(Lsu2Plugin_setup_sharedCompletion_valid) begin
      _zz_7 = 1'b1;
    end
  end

  always @(*) begin
    _zz_8 = 1'b0;
    if(RobPlugin_logic_completionMem_targetWrite_valid) begin
      _zz_8 = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid = 1'b0;
    if(BranchContextPlugin_free_dispatchMem_writes_1_port_valid) begin
      _zz_io_writes_1_valid = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_writes_0_valid = 1'b0;
    if(BranchContextPlugin_free_dispatchMem_writes_0_port_valid) begin
      _zz_io_writes_0_valid = 1'b1;
    end
  end

  always @(*) begin
    DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_2 = DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_1;
    if(when_DecoderPredictionPlugin_l212_1) begin
      DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_2 = 1'b1;
    end
  end

  always @(*) begin
    DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_1 = DecoderPredictionPlugin_logic_decodePatch_rasPushUsed;
    if(when_DecoderPredictionPlugin_l212) begin
      DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_9 = 1'b0;
    if(CsrRamPlugin_logic_writeLogic_port_valid) begin
      _zz_9 = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid_1 = 1'b0;
    if(ALU1_BranchPlugin_logic_branch_finalBranch_valid) begin
      _zz_io_writes_1_valid_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_writes_0_valid_1 = 1'b0;
    if(ALU0_BranchPlugin_logic_branch_finalBranch_valid) begin
      _zz_io_writes_0_valid_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548 = 1'b0;
    if(Lsu2Plugin_logic_flush_busy) begin
      _zz_FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548 = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_writes_2_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(!when_Lsu2Plugin_l1374) begin
              _zz_io_writes_2_valid = 1'b1;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    _zz_io_writes_2_valid_1 = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(!when_Lsu2Plugin_l1333) begin
              _zz_io_writes_2_valid_1 = 1'b1;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid_2 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_io_writes_1_valid_2 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_10 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_10 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_11 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_11 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid_3 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_io_writes_1_valid_3 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_12 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_12 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_13 = 1'b0;
    if(when_Lsu2Plugin_l1052) begin
      if(Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) begin
        _zz_13 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_2_valid_2 = 1'b0;
    if(when_Lsu2Plugin_l959) begin
      _zz_io_writes_2_valid_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842 = 1'b0;
    if(when_Lsu2Plugin_l841) begin
      _zz_Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842 = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_allocation_stores_alloc_2 = Lsu2Plugin_logic_allocation_stores_alloc_1;
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      Lsu2Plugin_logic_allocation_stores_alloc_2 = (Lsu2Plugin_logic_allocation_stores_alloc_1 + 5'h01);
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid_4 = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_1_valid_4 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid_5 = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_1_valid_5 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid_6 = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_1_valid_6 = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_allocation_loads_alloc_2 = Lsu2Plugin_logic_allocation_loads_alloc_1;
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      Lsu2Plugin_logic_allocation_loads_alloc_2 = (Lsu2Plugin_logic_allocation_loads_alloc_1 + 5'h01);
    end
  end

  always @(*) begin
    _zz_14 = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_14 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid_7 = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_1_valid_7 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid_8 = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_1_valid_8 = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_allocation_stores_alloc_1 = Lsu2Plugin_logic_allocation_stores_alloc;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      Lsu2Plugin_logic_allocation_stores_alloc_1 = (Lsu2Plugin_logic_allocation_stores_alloc + 5'h01);
    end
  end

  always @(*) begin
    _zz_io_writes_0_valid_2 = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_0_valid_2 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_0_valid_3 = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_0_valid_3 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_0_valid_4 = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_0_valid_4 = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_allocation_loads_alloc_1 = Lsu2Plugin_logic_allocation_loads_alloc;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      Lsu2Plugin_logic_allocation_loads_alloc_1 = (Lsu2Plugin_logic_allocation_loads_alloc + 5'h01);
    end
  end

  always @(*) begin
    _zz_15 = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_15 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_0_valid_5 = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_0_valid_5 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_io_writes_0_valid_6 = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        _zz_io_writes_0_valid_6 = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_onCommit_commitComb_2 = Lsu2Plugin_logic_sq_onCommit_commitComb_1;
    Lsu2Plugin_logic_sq_onCommit_commitComb_2 = (Lsu2Plugin_logic_sq_onCommit_commitComb_1 + _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_2);
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_onCommit_commitComb_1 = Lsu2Plugin_logic_sq_onCommit_commitComb;
    Lsu2Plugin_logic_sq_onCommit_commitComb_1 = (Lsu2Plugin_logic_sq_onCommit_commitComb + _zz_Lsu2Plugin_logic_sq_onCommit_commitComb_1);
  end

  always @(*) begin
    _zz_when_MultiportRam_l362 = 1'b0;
    if(Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_valid) begin
      _zz_when_MultiportRam_l362 = 1'b1;
    end
  end

  always @(*) begin
    _zz_when_MultiportRam_l362_1 = 1'b0;
    if(Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_valid) begin
      _zz_when_MultiportRam_l362_1 = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_onCommit_free_2 = Lsu2Plugin_logic_lq_onCommit_free_1;
    Lsu2Plugin_logic_lq_onCommit_free_2 = (Lsu2Plugin_logic_lq_onCommit_free_1 + _zz_Lsu2Plugin_logic_lq_onCommit_free_2);
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_onCommit_priority_2 = Lsu2Plugin_logic_lq_onCommit_priority_1;
    if(Lsu2Plugin_logic_lq_onCommit_lqCommits_1) begin
      Lsu2Plugin_logic_lq_onCommit_priority_2 = ((Lsu2Plugin_logic_lq_onCommit_priority_1 == 15'h0000) ? 15'h7fff : _zz_Lsu2Plugin_logic_lq_onCommit_priority_2);
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_onCommit_free_1 = Lsu2Plugin_logic_lq_onCommit_free;
    Lsu2Plugin_logic_lq_onCommit_free_1 = (Lsu2Plugin_logic_lq_onCommit_free + _zz_Lsu2Plugin_logic_lq_onCommit_free_1);
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_onCommit_priority_1 = Lsu2Plugin_logic_lq_onCommit_priority;
    if(Lsu2Plugin_logic_lq_onCommit_lqCommits_0) begin
      Lsu2Plugin_logic_lq_onCommit_priority_1 = ((Lsu2Plugin_logic_lq_onCommit_priority == 15'h0000) ? 15'h7fff : _zz_Lsu2Plugin_logic_lq_onCommit_priority_1);
    end
  end

  always @(*) begin
    HistoryPlugin_logic_update_pushes_2_stateNext_2 = HistoryPlugin_logic_update_pushes_2_stateNext_1;
    if(when_HistoryPlugin_l115_2) begin
      HistoryPlugin_logic_update_pushes_2_stateNext_2 = _zz_HistoryPlugin_logic_update_pushes_2_stateNext_2[23:0];
    end
  end

  always @(*) begin
    HistoryPlugin_logic_update_pushes_2_stateNext_1 = HistoryPlugin_logic_update_pushes_2_stateNext;
    if(when_HistoryPlugin_l115_1) begin
      HistoryPlugin_logic_update_pushes_2_stateNext_1 = _zz_HistoryPlugin_logic_update_pushes_2_stateNext_1[23:0];
    end
  end

  always @(*) begin
    HistoryPlugin_logic_update_pushes_0_stateNext_1 = HistoryPlugin_logic_update_pushes_0_stateNext;
    if(when_HistoryPlugin_l115) begin
      HistoryPlugin_logic_update_pushes_0_stateNext_1 = _zz_HistoryPlugin_logic_update_pushes_0_stateNext_1[23:0];
    end
  end

  always @(*) begin
    HistoryPlugin_logic_onCommit_valueNext_2 = HistoryPlugin_logic_onCommit_valueNext_1;
    if(when_HistoryPlugin_l90_1) begin
      HistoryPlugin_logic_onCommit_valueNext_2 = _zz_HistoryPlugin_logic_onCommit_valueNext_2[23:0];
    end
  end

  always @(*) begin
    HistoryPlugin_logic_onCommit_valueNext_1 = HistoryPlugin_logic_onCommit_valueNext;
    if(when_HistoryPlugin_l90) begin
      HistoryPlugin_logic_onCommit_valueNext_1 = _zz_HistoryPlugin_logic_onCommit_valueNext_1[23:0];
    end
  end

  always @(*) begin
    CommitPlugin_logic_commit_continue_2 = CommitPlugin_logic_commit_continue_1;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_commit_slot_1_enable) begin
        if(when_CommitPlugin_l211_1) begin
          CommitPlugin_logic_commit_continue_2 = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    CommitPlugin_logic_commit_continue_1 = CommitPlugin_logic_commit_continue;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_commit_slot_0_enable) begin
        if(when_CommitPlugin_l211) begin
          CommitPlugin_logic_commit_continue_1 = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    _zz_when_MultiportRam_l328 = 1'b0;
    if(GSharePlugin_logic_mem_write_valid) begin
      _zz_when_MultiportRam_l328 = 1'b1;
    end
  end

  always @(*) begin
    _zz_16 = 1'b0;
    if(BtbPlugin_logic_onLearn_port_valid) begin
      _zz_16 = 1'b1;
    end
  end

  always @(*) begin
    _zz_17 = 1'b0;
    if(DecoderPredictionPlugin_logic_ras_write_valid) begin
      _zz_17 = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid_9 = 1'b0;
    if(when_BranchContextPlugin_l93_1) begin
      if(FrontendPlugin_allocated_ready) begin
        _zz_io_writes_1_valid_9 = 1'b1;
      end
    end
  end

  always @(*) begin
    BranchContextPlugin_logic_alloc_allocNext_2 = BranchContextPlugin_logic_alloc_allocNext_1;
    if(when_BranchContextPlugin_l93_1) begin
      BranchContextPlugin_logic_alloc_allocNext_2 = (BranchContextPlugin_logic_alloc_allocNext_1 + 5'h01);
    end
  end

  always @(*) begin
    _zz_io_writes_0_valid_7 = 1'b0;
    if(when_BranchContextPlugin_l93) begin
      if(FrontendPlugin_allocated_ready) begin
        _zz_io_writes_0_valid_7 = 1'b1;
      end
    end
  end

  always @(*) begin
    BranchContextPlugin_logic_alloc_allocNext_1 = BranchContextPlugin_logic_alloc_allocNext;
    if(when_BranchContextPlugin_l93) begin
      BranchContextPlugin_logic_alloc_allocNext_1 = (BranchContextPlugin_logic_alloc_allocNext + 5'h01);
    end
  end

  always @(*) begin
    AlignerPlugin_logic_slices_remains_2 = AlignerPlugin_logic_slices_remains_1;
    AlignerPlugin_logic_slices_remains_2 = (AlignerPlugin_logic_slices_remains_1 & (~ (AlignerPlugin_logic_extractors_1_valid ? AlignerPlugin_logic_extractors_1_usage : 4'b0000)));
  end

  always @(*) begin
    AlignerPlugin_logic_slices_carry_2 = AlignerPlugin_logic_slices_carry_1;
    AlignerPlugin_logic_slices_carry_2 = (AlignerPlugin_logic_slices_carry_1 & (~ AlignerPlugin_logic_extractors_1_usage));
  end

  always @(*) begin
    AlignerPlugin_logic_slices_used_2 = AlignerPlugin_logic_slices_used_1;
    AlignerPlugin_logic_slices_used_2 = (AlignerPlugin_logic_slices_used_1 | AlignerPlugin_logic_extractors_1_usage);
  end

  always @(*) begin
    AlignerPlugin_logic_slices_remains_1 = AlignerPlugin_logic_slices_remains;
    AlignerPlugin_logic_slices_remains_1 = (AlignerPlugin_logic_slices_remains & (~ (AlignerPlugin_logic_extractors_0_valid ? AlignerPlugin_logic_extractors_0_usage : 4'b0000)));
  end

  always @(*) begin
    AlignerPlugin_logic_slices_carry_1 = AlignerPlugin_logic_slices_carry;
    AlignerPlugin_logic_slices_carry_1 = (AlignerPlugin_logic_slices_carry & (~ AlignerPlugin_logic_extractors_0_usage));
  end

  always @(*) begin
    AlignerPlugin_logic_slices_used_1 = AlignerPlugin_logic_slices_used;
    AlignerPlugin_logic_slices_used_1 = (AlignerPlugin_logic_slices_used | AlignerPlugin_logic_extractors_0_usage);
  end

  always @(*) begin
    _zz_FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552 = 1'b0;
    if(FetchCachePlugin_logic_read_ctrl_redoIt) begin
      _zz_FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552 = 1'b1;
    end
  end

  always @(*) begin
    _zz_FetchPlugin_stages_2_isFlushingRoot = 1'b0;
    if(FetchCachePlugin_logic_read_ctrl_redoIt) begin
      _zz_FetchPlugin_stages_2_isFlushingRoot = 1'b1;
    end
  end

  always @(*) begin
    _zz_18 = 1'b0;
    if(FetchCachePlugin_logic_plru_write_valid) begin
      _zz_18 = 1'b1;
    end
  end

  always @(*) begin
    _zz_when_MultiportRam_l328_1 = 1'b0;
    if(FetchCachePlugin_logic_banks_3_write_valid) begin
      _zz_when_MultiportRam_l328_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_when_MultiportRam_l328_2 = 1'b0;
    if(FetchCachePlugin_logic_banks_2_write_valid) begin
      _zz_when_MultiportRam_l328_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_when_MultiportRam_l328_3 = 1'b0;
    if(FetchCachePlugin_logic_banks_1_write_valid) begin
      _zz_when_MultiportRam_l328_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_when_MultiportRam_l328_4 = 1'b0;
    if(FetchCachePlugin_logic_banks_0_write_valid) begin
      _zz_when_MultiportRam_l328_4 = 1'b1;
    end
  end

  always @(*) begin
    PcPlugin_logic_jump_target_1 = PcPlugin_logic_jump_target;
    if(when_PcPlugin_l55) begin
      PcPlugin_logic_jump_target_1 = (_zz_PcPlugin_logic_jump_target_1 ? BtbPlugin_setup_btbJump_payload_pc : 32'h00000000);
    end
  end

  always @(*) begin
    MmuPlugin_setup_invalidatePort_cmd_valid = 1'b0;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
        if(EnvCallPlugin_logic_flushes_vmaInv) begin
          MmuPlugin_setup_invalidatePort_cmd_valid = 1'b1;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
    if(when_CsrAccessPlugin_l181) begin
      MmuPlugin_setup_invalidatePort_cmd_valid = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_setup_invalidatePort_rsp_valid = 1'b0;
    if(when_MmuPlugin_l515) begin
      MmuPlugin_setup_invalidatePort_rsp_valid = 1'b1;
    end
  end

  always @(*) begin
    FetchCachePlugin_setup_invalidatePort_cmd_valid = 1'b0;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
        if(EnvCallPlugin_logic_flushes_fetchInv) begin
          FetchCachePlugin_setup_invalidatePort_cmd_valid = 1'b1;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_invalidatePort_rsp_valid = 1'b0;
    if(when_FetchCachePlugin_l400) begin
      FetchCachePlugin_setup_invalidatePort_rsp_valid = 1'b1;
    end
  end

  assign AlignerPlugin_setup_singleFetch = 1'b0;
  assign FrontendPlugin_decoded_isFireing = (FrontendPlugin_decoded_valid && FrontendPlugin_decoded_ready);
  assign FrontendPlugin_allocated_isFireing = (FrontendPlugin_allocated_valid && FrontendPlugin_allocated_ready);
  always @(*) begin
    DecoderPlugin_setup_trapHalt = 1'b0;
    if(PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt) begin
      DecoderPlugin_setup_trapHalt = 1'b1;
    end
  end

  always @(*) begin
    DecoderPlugin_setup_trapRaise = 1'b0;
    if(when_PrivilegedPlugin_l672) begin
      DecoderPlugin_setup_trapRaise = 1'b1;
    end
  end

  assign DecoderPlugin_setup_debugEnter_0 = 1'b0;
  assign DecoderPlugin_setup_debugEnter_1 = 1'b0;
  always @(*) begin
    Lsu2Plugin_setup_postCommitBusy = 1'b0;
    if(when_Lsu2Plugin_l572) begin
      Lsu2Plugin_setup_postCommitBusy = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_flushPort_cmd_valid = 1'b0;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
        Lsu2Plugin_setup_flushPort_cmd_valid = 1'b1;
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_flushPort_cmd_payload_withFree = 1'bx;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
        Lsu2Plugin_setup_flushPort_cmd_payload_withFree = EnvCallPlugin_logic_flushes_flushData;
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_flushPort_rsp_valid = 1'b0;
    if(when_Lsu2Plugin_l1553) begin
      if(when_Lsu2Plugin_l1569) begin
        Lsu2Plugin_setup_flushPort_rsp_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    PrivilegedPlugin_setup_jump_valid = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
        PrivilegedPlugin_setup_jump_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
        PrivilegedPlugin_setup_jump_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_setup_jump_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_jump_payload_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
        PrivilegedPlugin_setup_jump_payload_pc = PrivilegedPlugin_logic_readed;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
        PrivilegedPlugin_setup_jump_payload_pc = PrivilegedPlugin_logic_readed;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_setup_jump_payload_pc = PrivilegedPlugin_logic_readed;
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_setup_withMachinePrivilege = (2'b11 <= PrivilegedPlugin_setup_privilege);
  assign PrivilegedPlugin_setup_withSupervisorPrivilege = (2'b01 <= PrivilegedPlugin_setup_privilege);
  always @(*) begin
    PrivilegedPlugin_setup_xretAwayFromMachine = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
        if(when_PrivilegedPlugin_l952) begin
          PrivilegedPlugin_setup_xretAwayFromMachine = 1'b1;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_trapEvent = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_setup_trapEvent = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_redoTriggered = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
        if(!when_PrivilegedPlugin_l766) begin
          case(PrivilegedPlugin_logic_reschedule_payload_cause)
            4'b1001 : begin
            end
            4'b1010 : begin
              PrivilegedPlugin_setup_redoTriggered = 1'b1;
            end
            4'b1000 : begin
            end
            default : begin
            end
          endcase
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_setup_setFpDirty = 1'b0;
  assign PrivilegedPlugin_setup_isFpuEnabled = 1'b0;
  always @(*) begin
    EU0_CsrAccessPlugin_setup_onDecodeTrap = 1'b0;
    if(when_PrivilegedPlugin_l165) begin
      EU0_CsrAccessPlugin_setup_onDecodeTrap = 1'b1;
    end
    if(when_PerformanceCounterPlugin_l268) begin
      EU0_CsrAccessPlugin_setup_onDecodeTrap = 1'b1;
    end
  end

  always @(*) begin
    EU0_CsrAccessPlugin_setup_onDecodeFlushPipeline = 1'b0;
    if(when_CsrAccessPlugin_l181) begin
      EU0_CsrAccessPlugin_setup_onDecodeFlushPipeline = 1'b1;
    end
  end

  always @(*) begin
    EU0_CsrAccessPlugin_setup_onReadHalt = 1'b0;
    if(PerformanceCounterPlugin_logic_csrRead_requested) begin
      if(when_PerformanceCounterPlugin_l253) begin
        EU0_CsrAccessPlugin_setup_onReadHalt = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l270) begin
      EU0_CsrAccessPlugin_setup_onReadHalt = 1'b1;
    end
  end

  always @(*) begin
    EU0_CsrAccessPlugin_setup_onWriteHalt = 1'b0;
    if(when_CsrAccessPlugin_l325) begin
      if(when_PerformanceCounterPlugin_l273) begin
        if(when_PerformanceCounterPlugin_l275) begin
          EU0_CsrAccessPlugin_setup_onWriteHalt = 1'b1;
        end
      end
    end
    if(when_CsrAccessPlugin_l340) begin
      EU0_CsrAccessPlugin_setup_onWriteHalt = 1'b1;
    end
  end

  assign EU0_CsrAccessPlugin_setup_onWriteFlushPipeline = 1'b0;
  assign FetchPlugin_stages_1_isFireing = (FetchPlugin_stages_1_valid && FetchPlugin_stages_1_ready);
  assign when_Stage_l170 = (FetchPlugin_stages_1_ready || FetchPlugin_stages_1_isFlushed);
  assign FetchPlugin_stages_1_isFirstCycle = (FetchPlugin_stages_1_valid && (! _zz_FetchPlugin_stages_1_isFirstCycle));
  assign _zz_PcPlugin_logic_jump_oh = {BtbPlugin_setup_btbJump_valid,{FetchCachePlugin_setup_redoJump_valid,{AlignerPlugin_setup_sequenceJump_valid,{DecoderPredictionPlugin_setup_decodeJump_valid,{CommitPlugin_setup_jump_valid,PrivilegedPlugin_setup_jump_valid}}}}};
  assign _zz_PcPlugin_logic_jump_oh_1 = _zz_PcPlugin_logic_jump_oh[0];
  assign _zz_PcPlugin_logic_jump_oh_2 = _zz_PcPlugin_logic_jump_oh[1];
  assign _zz_PcPlugin_logic_jump_oh_3 = _zz_PcPlugin_logic_jump_oh[2];
  assign _zz_PcPlugin_logic_jump_oh_4 = _zz_PcPlugin_logic_jump_oh[3];
  assign _zz_PcPlugin_logic_jump_oh_5 = _zz_PcPlugin_logic_jump_oh[4];
  always @(*) begin
    _zz_PcPlugin_logic_jump_oh_6[0] = (_zz_PcPlugin_logic_jump_oh_1 && (! 1'b0));
    _zz_PcPlugin_logic_jump_oh_6[1] = (_zz_PcPlugin_logic_jump_oh_2 && (! _zz_PcPlugin_logic_jump_oh_1));
    _zz_PcPlugin_logic_jump_oh_6[2] = (_zz_PcPlugin_logic_jump_oh_3 && (! ({_zz_PcPlugin_logic_jump_oh_2,_zz_PcPlugin_logic_jump_oh_1} != 2'b00)));
    _zz_PcPlugin_logic_jump_oh_6[3] = (_zz_PcPlugin_logic_jump_oh_4 && (! ({_zz_PcPlugin_logic_jump_oh_3,{_zz_PcPlugin_logic_jump_oh_2,_zz_PcPlugin_logic_jump_oh_1}} != 3'b000)));
    _zz_PcPlugin_logic_jump_oh_6[4] = (_zz_PcPlugin_logic_jump_oh_5 && (! ({_zz_PcPlugin_logic_jump_oh_4,{_zz_PcPlugin_logic_jump_oh_3,{_zz_PcPlugin_logic_jump_oh_2,_zz_PcPlugin_logic_jump_oh_1}}} != 4'b0000)));
    _zz_PcPlugin_logic_jump_oh_6[5] = (_zz_PcPlugin_logic_jump_oh[5] && (! ({_zz_PcPlugin_logic_jump_oh_5,{_zz_PcPlugin_logic_jump_oh_4,{_zz_PcPlugin_logic_jump_oh_3,{_zz_PcPlugin_logic_jump_oh_2,_zz_PcPlugin_logic_jump_oh_1}}}} != 5'h00)));
  end

  assign PcPlugin_logic_jump_oh = _zz_PcPlugin_logic_jump_oh_6;
  assign PcPlugin_logic_jump_target = ((((PcPlugin_logic_jump_oh[0] ? PrivilegedPlugin_setup_jump_payload_pc : 32'h00000000) | (PcPlugin_logic_jump_oh[1] ? CommitPlugin_setup_jump_payload_pc : 32'h00000000)) | ((PcPlugin_logic_jump_oh[2] ? DecoderPredictionPlugin_setup_decodeJump_payload_pc : 32'h00000000) | (PcPlugin_logic_jump_oh[3] ? AlignerPlugin_setup_sequenceJump_payload_pc : 32'h00000000))) | (PcPlugin_logic_jump_oh[4] ? FetchCachePlugin_setup_redoJump_payload_pc : 32'h00000000));
  assign _zz_PcPlugin_logic_jump_target_1 = PcPlugin_logic_jump_oh[5];
  assign when_PcPlugin_l55 = (_zz_PcPlugin_logic_jump_target_1 != 1'b0);
  assign PcPlugin_logic_jump_pcLoad_valid = ({PrivilegedPlugin_setup_jump_valid,{CommitPlugin_setup_jump_valid,{BtbPlugin_setup_btbJump_valid,{DecoderPredictionPlugin_setup_decodeJump_valid,{AlignerPlugin_setup_sequenceJump_valid,FetchCachePlugin_setup_redoJump_valid}}}}} != 6'h00);
  assign PcPlugin_logic_jump_pcLoad_payload_pc = PcPlugin_logic_jump_target_1;
  assign FetchCachePlugin_logic_banks_0_read_rsp = _zz_FetchCachePlugin_logic_banks_0_read_rsp;
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_0 = FetchCachePlugin_logic_banks_0_read_rsp;
  assign FetchCachePlugin_logic_banks_1_read_rsp = _zz_FetchCachePlugin_logic_banks_1_read_rsp;
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_1 = FetchCachePlugin_logic_banks_1_read_rsp;
  assign FetchCachePlugin_logic_banks_2_read_rsp = _zz_FetchCachePlugin_logic_banks_2_read_rsp;
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_2 = FetchCachePlugin_logic_banks_2_read_rsp;
  assign FetchCachePlugin_logic_banks_3_read_rsp = _zz_FetchCachePlugin_logic_banks_3_read_rsp;
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_3 = FetchCachePlugin_logic_banks_3_read_rsp;
  always @(*) begin
    FetchCachePlugin_logic_waysWrite_mask = 4'b0000;
    if(when_FetchCachePlugin_l383) begin
      FetchCachePlugin_logic_waysWrite_mask = 4'b1111;
    end
    if(FetchCachePlugin_logic_invalidate_done) begin
      if(FetchCachePlugin_logic_refill_fire) begin
        FetchCachePlugin_logic_waysWrite_mask[FetchCachePlugin_logic_refill_wayToAllocate] = 1'b1;
      end
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_waysWrite_address = 6'bxxxxxx;
    if(when_FetchCachePlugin_l383) begin
      FetchCachePlugin_logic_waysWrite_address = FetchCachePlugin_logic_invalidate_counter[5:0];
    end
    if(FetchCachePlugin_logic_invalidate_done) begin
      FetchCachePlugin_logic_waysWrite_address = FetchCachePlugin_logic_refill_address[11 : 6];
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_waysWrite_tag_loaded = 1'bx;
    if(when_FetchCachePlugin_l383) begin
      FetchCachePlugin_logic_waysWrite_tag_loaded = 1'b0;
    end
    if(FetchCachePlugin_logic_invalidate_done) begin
      FetchCachePlugin_logic_waysWrite_tag_loaded = 1'b1;
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_waysWrite_tag_error = 1'bx;
    if(FetchCachePlugin_logic_invalidate_done) begin
      FetchCachePlugin_logic_waysWrite_tag_error = (FetchCachePlugin_logic_refill_hadError || FetchCachePlugin_mem_rsp_payload_error);
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(FetchCachePlugin_logic_invalidate_done) begin
      FetchCachePlugin_logic_waysWrite_tag_address = FetchCachePlugin_logic_refill_address[31 : 12];
    end
  end

  assign _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded = _zz_FetchCachePlugin_logic_ways_0_mem_port1;
  assign FetchCachePlugin_logic_ways_0_read_rsp_loaded = _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded[0];
  assign FetchCachePlugin_logic_ways_0_read_rsp_error = _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded[1];
  assign FetchCachePlugin_logic_ways_0_read_rsp_address = _zz_FetchCachePlugin_logic_ways_0_read_rsp_loaded[21 : 2];
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_loaded = FetchCachePlugin_logic_ways_0_read_rsp_loaded;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_error = FetchCachePlugin_logic_ways_0_read_rsp_error;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_address = FetchCachePlugin_logic_ways_0_read_rsp_address;
  assign _zz_FetchCachePlugin_logic_ways_1_read_rsp_loaded = _zz_FetchCachePlugin_logic_ways_1_mem_port1;
  assign FetchCachePlugin_logic_ways_1_read_rsp_loaded = _zz_FetchCachePlugin_logic_ways_1_read_rsp_loaded[0];
  assign FetchCachePlugin_logic_ways_1_read_rsp_error = _zz_FetchCachePlugin_logic_ways_1_read_rsp_loaded[1];
  assign FetchCachePlugin_logic_ways_1_read_rsp_address = _zz_FetchCachePlugin_logic_ways_1_read_rsp_loaded[21 : 2];
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_1_loaded = FetchCachePlugin_logic_ways_1_read_rsp_loaded;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_1_error = FetchCachePlugin_logic_ways_1_read_rsp_error;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_1_address = FetchCachePlugin_logic_ways_1_read_rsp_address;
  assign _zz_FetchCachePlugin_logic_ways_2_read_rsp_loaded = _zz_FetchCachePlugin_logic_ways_2_mem_port1;
  assign FetchCachePlugin_logic_ways_2_read_rsp_loaded = _zz_FetchCachePlugin_logic_ways_2_read_rsp_loaded[0];
  assign FetchCachePlugin_logic_ways_2_read_rsp_error = _zz_FetchCachePlugin_logic_ways_2_read_rsp_loaded[1];
  assign FetchCachePlugin_logic_ways_2_read_rsp_address = _zz_FetchCachePlugin_logic_ways_2_read_rsp_loaded[21 : 2];
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_2_loaded = FetchCachePlugin_logic_ways_2_read_rsp_loaded;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_2_error = FetchCachePlugin_logic_ways_2_read_rsp_error;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_2_address = FetchCachePlugin_logic_ways_2_read_rsp_address;
  assign _zz_FetchCachePlugin_logic_ways_3_read_rsp_loaded = _zz_FetchCachePlugin_logic_ways_3_mem_port1;
  assign FetchCachePlugin_logic_ways_3_read_rsp_loaded = _zz_FetchCachePlugin_logic_ways_3_read_rsp_loaded[0];
  assign FetchCachePlugin_logic_ways_3_read_rsp_error = _zz_FetchCachePlugin_logic_ways_3_read_rsp_loaded[1];
  assign FetchCachePlugin_logic_ways_3_read_rsp_address = _zz_FetchCachePlugin_logic_ways_3_read_rsp_loaded[21 : 2];
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_3_loaded = FetchCachePlugin_logic_ways_3_read_rsp_loaded;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_3_error = FetchCachePlugin_logic_ways_3_read_rsp_error;
  assign FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_3_address = FetchCachePlugin_logic_ways_3_read_rsp_address;
  always @(*) begin
    FetchCachePlugin_logic_invalidate_canStart = 1'b1;
    if(when_FetchCachePlugin_l396) begin
      FetchCachePlugin_logic_invalidate_canStart = 1'b0;
    end
    if(FetchCachePlugin_logic_refill_valid) begin
      FetchCachePlugin_logic_invalidate_canStart = 1'b0;
    end
  end

  assign FetchCachePlugin_logic_invalidate_done = FetchCachePlugin_logic_invalidate_counter[6];
  assign when_FetchCachePlugin_l379 = (! FetchCachePlugin_logic_invalidate_done);
  assign when_FetchCachePlugin_l383 = (! FetchCachePlugin_logic_invalidate_done);
  assign FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l389 = ((! FetchCachePlugin_logic_invalidate_done) || FetchCachePlugin_logic_invalidate_requested);
  assign when_FetchCachePlugin_l391 = (FetchCachePlugin_logic_invalidate_requested && FetchCachePlugin_logic_invalidate_canStart);
  assign when_FetchCachePlugin_l396 = ({FetchPlugin_stages_2_valid,FetchPlugin_stages_1_valid} != 2'b00);
  assign when_FetchCachePlugin_l400 = (FetchCachePlugin_logic_invalidate_done && (! FetchCachePlugin_logic_invalidate_done_regNext));
  always @(*) begin
    FetchCachePlugin_logic_refill_start_valid = 1'b0;
    if(FetchPlugin_stages_2_valid) begin
      if(!FetchPlugin_stages_2_MMU_REDO) begin
        if(when_FetchCachePlugin_l562) begin
          FetchCachePlugin_logic_refill_start_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_refill_fire = 1'b0;
    if(FetchCachePlugin_mem_rsp_valid) begin
      if(when_FetchCachePlugin_l470) begin
        FetchCachePlugin_logic_refill_fire = 1'b1;
      end
    end
  end

  assign when_FetchCachePlugin_l422 = (! FetchCachePlugin_logic_refill_valid);
  assign FetchCachePlugin_mem_cmd_fire = (FetchCachePlugin_mem_cmd_valid && FetchCachePlugin_mem_cmd_ready);
  assign FetchCachePlugin_mem_cmd_valid = (FetchCachePlugin_logic_refill_valid && (! FetchCachePlugin_logic_refill_cmdSent));
  assign FetchCachePlugin_mem_cmd_payload_address = {FetchCachePlugin_logic_refill_address[31 : 6],6'h00};
  assign FetchCachePlugin_mem_cmd_payload_io = FetchCachePlugin_logic_refill_isIo;
  assign when_Utils_l560 = (! FetchCachePlugin_logic_refill_valid);
  always @(*) begin
    FetchCachePlugin_logic_refill_randomWay_willIncrement = 1'b0;
    if(when_Utils_l560) begin
      FetchCachePlugin_logic_refill_randomWay_willIncrement = 1'b1;
    end
  end

  assign FetchCachePlugin_logic_refill_randomWay_willClear = 1'b0;
  assign FetchCachePlugin_logic_refill_randomWay_willOverflowIfInc = (FetchCachePlugin_logic_refill_randomWay_value == 2'b11);
  assign FetchCachePlugin_logic_refill_randomWay_willOverflow = (FetchCachePlugin_logic_refill_randomWay_willOverflowIfInc && FetchCachePlugin_logic_refill_randomWay_willIncrement);
  always @(*) begin
    FetchCachePlugin_logic_refill_randomWay_valueNext = (FetchCachePlugin_logic_refill_randomWay_value + _zz_FetchCachePlugin_logic_refill_randomWay_valueNext);
    if(FetchCachePlugin_logic_refill_randomWay_willClear) begin
      FetchCachePlugin_logic_refill_randomWay_valueNext = 2'b00;
    end
  end

  assign FetchCachePlugin_logic_banks_0_write_valid = (FetchCachePlugin_mem_rsp_valid && (FetchCachePlugin_logic_refill_wayToAllocate == 2'b00));
  assign FetchCachePlugin_logic_banks_0_write_payload_address = {FetchCachePlugin_logic_refill_address[11 : 6],FetchCachePlugin_logic_refill_wordIndex};
  assign FetchCachePlugin_logic_banks_0_write_payload_data = FetchCachePlugin_mem_rsp_payload_data;
  assign FetchCachePlugin_logic_banks_1_write_valid = (FetchCachePlugin_mem_rsp_valid && (FetchCachePlugin_logic_refill_wayToAllocate == 2'b01));
  assign FetchCachePlugin_logic_banks_1_write_payload_address = {FetchCachePlugin_logic_refill_address[11 : 6],FetchCachePlugin_logic_refill_wordIndex};
  assign FetchCachePlugin_logic_banks_1_write_payload_data = FetchCachePlugin_mem_rsp_payload_data;
  assign FetchCachePlugin_logic_banks_2_write_valid = (FetchCachePlugin_mem_rsp_valid && (FetchCachePlugin_logic_refill_wayToAllocate == 2'b10));
  assign FetchCachePlugin_logic_banks_2_write_payload_address = {FetchCachePlugin_logic_refill_address[11 : 6],FetchCachePlugin_logic_refill_wordIndex};
  assign FetchCachePlugin_logic_banks_2_write_payload_data = FetchCachePlugin_mem_rsp_payload_data;
  assign FetchCachePlugin_logic_banks_3_write_valid = (FetchCachePlugin_mem_rsp_valid && (FetchCachePlugin_logic_refill_wayToAllocate == 2'b11));
  assign FetchCachePlugin_logic_banks_3_write_payload_address = {FetchCachePlugin_logic_refill_address[11 : 6],FetchCachePlugin_logic_refill_wordIndex};
  assign FetchCachePlugin_logic_banks_3_write_payload_data = FetchCachePlugin_mem_rsp_payload_data;
  assign FetchCachePlugin_mem_rsp_ready = 1'b1;
  assign when_FetchCachePlugin_l470 = (FetchCachePlugin_logic_refill_wordIndex == 3'b111);
  assign FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l476 = FetchCachePlugin_logic_refill_valid;
  assign FetchCachePlugin_setup_refillEvent = FetchCachePlugin_logic_refill_fire_regNext;
  assign FetchCachePlugin_logic_banks_0_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_banks_0_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[11 : 3];
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_0 = FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_0[63 : 0];
  assign FetchCachePlugin_logic_banks_1_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_banks_1_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[11 : 3];
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_1 = FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_1[63 : 0];
  assign FetchCachePlugin_logic_banks_2_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_banks_2_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[11 : 3];
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_2 = FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_2[63 : 0];
  assign FetchCachePlugin_logic_banks_3_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_banks_3_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[11 : 3];
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_3 = FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_WORDS_3[63 : 0];
  assign FetchPlugin_stages_2_Fetch_WORD = (((FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_0 ? FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_0 : 64'h0000000000000000) | (FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_1 ? FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_1 : 64'h0000000000000000)) | ((FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_2 ? FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_2 : 64'h0000000000000000) | (FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_3 ? FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_3 : 64'h0000000000000000)));
  assign FetchCachePlugin_logic_ways_0_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_ways_0_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[11 : 6];
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_0 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_0[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[0]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_1 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_1[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[1]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_2 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_2[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[2]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_3 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_3[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[3]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_4 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_4[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[4]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_5 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_5[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[5]);
  assign FetchCachePlugin_logic_read_onWays_0_hits_translatedHits = ({FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_5,{FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_4,{FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_3,{FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_2,{FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_1,FetchCachePlugin_logic_read_onWays_0_hits_wayTlbHits_0}}}}} != 6'h00);
  assign FetchCachePlugin_logic_read_onWays_0_hits_bypassHits = (FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address == _zz_FetchCachePlugin_logic_read_onWays_0_hits_bypassHits);
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_0 = ((FetchPlugin_stages_1_MMU_BYPASS_TRANSLATION ? FetchCachePlugin_logic_read_onWays_0_hits_bypassHits : FetchCachePlugin_logic_read_onWays_0_hits_translatedHits) && FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_loaded);
  assign FetchCachePlugin_logic_ways_1_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_ways_1_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[11 : 6];
  assign FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_0 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_0[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[0]);
  assign FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_1 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_1[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[1]);
  assign FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_2 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_2[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[2]);
  assign FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_3 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_3[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[3]);
  assign FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_4 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_4[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[4]);
  assign FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_5 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_5[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[5]);
  assign FetchCachePlugin_logic_read_onWays_1_hits_translatedHits = ({FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_5,{FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_4,{FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_3,{FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_2,{FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_1,FetchCachePlugin_logic_read_onWays_1_hits_wayTlbHits_0}}}}} != 6'h00);
  assign FetchCachePlugin_logic_read_onWays_1_hits_bypassHits = (FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address == _zz_FetchCachePlugin_logic_read_onWays_1_hits_bypassHits);
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_1 = ((FetchPlugin_stages_1_MMU_BYPASS_TRANSLATION ? FetchCachePlugin_logic_read_onWays_1_hits_bypassHits : FetchCachePlugin_logic_read_onWays_1_hits_translatedHits) && FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_loaded);
  assign FetchCachePlugin_logic_ways_2_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_ways_2_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[11 : 6];
  assign FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_0 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_0[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[0]);
  assign FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_1 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_1[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[1]);
  assign FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_2 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_2[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[2]);
  assign FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_3 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_3[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[3]);
  assign FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_4 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_4[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[4]);
  assign FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_5 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_5[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[5]);
  assign FetchCachePlugin_logic_read_onWays_2_hits_translatedHits = ({FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_5,{FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_4,{FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_3,{FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_2,{FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_1,FetchCachePlugin_logic_read_onWays_2_hits_wayTlbHits_0}}}}} != 6'h00);
  assign FetchCachePlugin_logic_read_onWays_2_hits_bypassHits = (FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address == _zz_FetchCachePlugin_logic_read_onWays_2_hits_bypassHits);
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_2 = ((FetchPlugin_stages_1_MMU_BYPASS_TRANSLATION ? FetchCachePlugin_logic_read_onWays_2_hits_bypassHits : FetchCachePlugin_logic_read_onWays_2_hits_translatedHits) && FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_loaded);
  assign FetchCachePlugin_logic_ways_3_read_cmd_valid = (! (FetchPlugin_stages_0_valid && (! FetchPlugin_stages_0_ready)));
  assign FetchCachePlugin_logic_ways_3_read_cmd_payload = FetchPlugin_stages_0_Fetch_FETCH_PC[11 : 6];
  assign FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_0 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_0[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[0]);
  assign FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_1 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_1[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[1]);
  assign FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_2 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_2[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[2]);
  assign FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_3 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_3[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[3]);
  assign FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_4 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_4[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[4]);
  assign FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_5 = ((FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address == FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_5[31 : 12]) && FetchPlugin_stages_1_MMU_WAYS_OH[5]);
  assign FetchCachePlugin_logic_read_onWays_3_hits_translatedHits = ({FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_5,{FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_4,{FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_3,{FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_2,{FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_1,FetchCachePlugin_logic_read_onWays_3_hits_wayTlbHits_0}}}}} != 6'h00);
  assign FetchCachePlugin_logic_read_onWays_3_hits_bypassHits = (FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address == _zz_FetchCachePlugin_logic_read_onWays_3_hits_bypassHits);
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_3 = ((FetchPlugin_stages_1_MMU_BYPASS_TRANSLATION ? FetchCachePlugin_logic_read_onWays_3_hits_bypassHits : FetchCachePlugin_logic_read_onWays_3_hits_translatedHits) && FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_loaded);
  assign _zz_FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0 = FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 6];
  assign _zz_FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0_1 = _zz_FetchCachePlugin_logic_plru_ram_port1;
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0 = _zz_FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0_1[0 : 0];
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_1 = _zz_FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0_1[2 : 1];
  assign FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HIT = (|{FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_3,{FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_2,{FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_1,FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_0}}});
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_logic_0_state = FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_context_state_0[0];
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_sel_0 = (! FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_logic_0_state);
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_logic_1_stateSel = FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_sel_0;
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_logic_1_state = FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_context_state_1[FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_logic_1_stateSel];
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_sel_1 = (! FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_logic_1_state);
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_evict_id = {FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_sel_0,FetchCachePlugin_logic_read_ctrl_plruLogic_core_evict_sel_1};
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_state_0[0] = FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id[1];
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_update_logic_1_sel = FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id[1 : 1];
  always @(*) begin
    FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_state_1 = FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_context_state_1;
    FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_state_1[FetchCachePlugin_logic_read_ctrl_plruLogic_core_update_logic_1_sel] = FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id[0];
  end

  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_context_state_0 = FetchPlugin_stages_2_FetchCachePlugin_logic_PLRU_0;
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_context_state_1 = FetchPlugin_stages_2_FetchCachePlugin_logic_PLRU_1;
  assign _zz_FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id = (FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_1 || FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_3);
  assign _zz_FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id_1 = (FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_2 || FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_3);
  assign FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id = {_zz_FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id_1,_zz_FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_id};
  always @(*) begin
    FetchCachePlugin_logic_plru_write_valid = 1'b0;
    if(!FetchCachePlugin_logic_read_ctrl_redoIt) begin
      if(FetchPlugin_stages_2_isFireing) begin
        FetchCachePlugin_logic_plru_write_valid = 1'b1;
      end
    end
    if(when_FetchCachePlugin_l593) begin
      FetchCachePlugin_logic_plru_write_valid = 1'b1;
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_plru_write_payload_address = FetchPlugin_stages_2_Fetch_FETCH_PC[11 : 6];
    if(when_FetchCachePlugin_l593) begin
      FetchCachePlugin_logic_plru_write_payload_address = FetchCachePlugin_logic_invalidate_counter[5:0];
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_plru_write_payload_data_0 = FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_state_0;
    if(when_FetchCachePlugin_l593) begin
      FetchCachePlugin_logic_plru_write_payload_data_0 = _zz_FetchCachePlugin_logic_plru_write_payload_data_0[0 : 0];
    end
  end

  always @(*) begin
    FetchCachePlugin_logic_plru_write_payload_data_1 = FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_update_state_1;
    if(when_FetchCachePlugin_l593) begin
      FetchCachePlugin_logic_plru_write_payload_data_1 = _zz_FetchCachePlugin_logic_plru_write_payload_data_0[2 : 1];
    end
  end

  assign FetchCachePlugin_logic_refill_start_wayToAllocate = FetchCachePlugin_logic_read_ctrl_plruLogic_core_io_evict_id;
  always @(*) begin
    FetchCachePlugin_setup_redoJump_valid = 1'b0;
    if(FetchCachePlugin_logic_read_ctrl_redoIt) begin
      FetchCachePlugin_setup_redoJump_valid = 1'b1;
    end
  end

  assign FetchCachePlugin_setup_redoJump_payload_pc = FetchPlugin_stages_2_Fetch_FETCH_PC;
  assign FetchPlugin_stages_2_Fetch_WORD_FAULT = (((|({FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_3,{FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_2,{FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_1,FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_0}}} & {FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_3_error,{FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_2_error,{FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_1_error,FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_error}}})) || FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE) || FetchPlugin_stages_2_MMU_ACCESS_FAULT);
  assign FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE = (FetchPlugin_stages_2_MMU_PAGE_FAULT || (! FetchPlugin_stages_2_MMU_ALLOW_EXECUTE));
  always @(*) begin
    FetchCachePlugin_logic_read_ctrl_redoIt = 1'b0;
    if(FetchPlugin_stages_2_valid) begin
      if(FetchPlugin_stages_2_MMU_REDO) begin
        FetchCachePlugin_logic_read_ctrl_redoIt = 1'b1;
      end else begin
        if(when_FetchCachePlugin_l562) begin
          FetchCachePlugin_logic_read_ctrl_redoIt = 1'b1;
        end
      end
    end
  end

  assign FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552 = _zz_FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552;
  assign FetchPlugin_stages_2_isFireing = (FetchPlugin_stages_2_valid && FetchPlugin_stages_2_ready);
  assign when_FetchCachePlugin_l562 = (((! FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE) && (! FetchPlugin_stages_2_MMU_ACCESS_FAULT)) && (! FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HIT));
  assign FetchCachePlugin_logic_refill_start_address = FetchPlugin_stages_2_MMU_TRANSLATED;
  assign FetchCachePlugin_logic_refill_start_isIo = FetchPlugin_stages_2_MMU_IO;
  assign FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l583 = (! FetchCachePlugin_logic_translationPort_wake);
  assign FetchCachePlugin_setup_historyJump_valid = FetchCachePlugin_setup_redoJump_valid;
  assign FetchCachePlugin_setup_historyJump_payload_history = FetchPlugin_stages_2_BRANCH_HISTORY;
  assign when_FetchCachePlugin_l593 = ((! FetchCachePlugin_logic_invalidate_done) && FetchCachePlugin_logic_invalidate_firstEver);
  assign _zz_FetchCachePlugin_logic_plru_write_payload_data_0 = 3'b000;
  assign AlignerPlugin_logic_ignoreInput = AlignerPlugin_setup_s2m_isFlushingRoot;
  assign AlignerPlugin_logic_isInputValid = (AlignerPlugin_setup_s2m_valid && (! AlignerPlugin_logic_ignoreInput));
  assign FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT = _zz_FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT;
  always @(*) begin
    AlignerPlugin_setup_s2m_MASK_BACK = _zz_AlignerPlugin_setup_s2m_MASK_BACK;
    if(when_AlignerPlugin_l98) begin
      AlignerPlugin_setup_s2m_MASK_BACK = 2'b11;
    end
  end

  assign when_AlignerPlugin_l98 = (! AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID);
  assign _zz_AlignerPlugin_logic_slices_data_0 = {AlignerPlugin_setup_s2m_Fetch_WORD,AlignerPlugin_logic_buffer_data};
  assign AlignerPlugin_logic_slices_data_0 = _zz_AlignerPlugin_logic_slices_data_0[31 : 0];
  assign AlignerPlugin_logic_slices_data_1 = _zz_AlignerPlugin_logic_slices_data_0[63 : 32];
  assign AlignerPlugin_logic_slices_data_2 = _zz_AlignerPlugin_logic_slices_data_0[95 : 64];
  assign AlignerPlugin_logic_slices_data_3 = _zz_AlignerPlugin_logic_slices_data_0[127 : 96];
  assign AlignerPlugin_logic_slices_carry = {(AlignerPlugin_logic_isInputValid ? AlignerPlugin_setup_s2m_MASK_FRONT : 2'b00),AlignerPlugin_logic_buffer_mask};
  assign AlignerPlugin_logic_slices_remains = AlignerPlugin_logic_slices_carry;
  assign AlignerPlugin_logic_slices_used = 4'b0000;
  assign AlignerPlugin_logic_decoders_0_usage = 4'b0001;
  assign AlignerPlugin_logic_decoders_0_notEnoughData = 1'b0;
  assign AlignerPlugin_logic_decoders_0_pastPrediction = 1'b0;
  assign AlignerPlugin_logic_decoders_0_usable = ((! AlignerPlugin_logic_decoders_0_notEnoughData) && (! AlignerPlugin_logic_decoders_0_pastPrediction));
  assign AlignerPlugin_logic_decoders_1_usage = 4'b0010;
  assign AlignerPlugin_logic_decoders_1_notEnoughData = 1'b0;
  assign AlignerPlugin_logic_decoders_1_pastPrediction = 1'b0;
  assign AlignerPlugin_logic_decoders_1_usable = ((! AlignerPlugin_logic_decoders_1_notEnoughData) && (! AlignerPlugin_logic_decoders_1_pastPrediction));
  assign AlignerPlugin_logic_decoders_2_usage = 4'b0100;
  assign AlignerPlugin_logic_decoders_2_notEnoughData = 1'b0;
  assign AlignerPlugin_logic_decoders_2_pastPrediction = 1'b0;
  assign AlignerPlugin_logic_decoders_2_usable = ((! AlignerPlugin_logic_decoders_2_notEnoughData) && (! AlignerPlugin_logic_decoders_2_pastPrediction));
  assign AlignerPlugin_logic_decoders_3_usage = 4'b1000;
  assign AlignerPlugin_logic_decoders_3_notEnoughData = 1'b0;
  assign AlignerPlugin_logic_decoders_3_pastPrediction = (AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID && (AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_SLICE < 1'b1));
  assign AlignerPlugin_logic_decoders_3_usable = ((! AlignerPlugin_logic_decoders_3_notEnoughData) && (! AlignerPlugin_logic_decoders_3_pastPrediction));
  assign _zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1 = 1'b0;
  assign _zz_AlignerPlugin_logic_extractors_0_maskOh = AlignerPlugin_logic_slices_carry[3 : 0];
  assign _zz_AlignerPlugin_logic_extractors_0_maskOh_1 = _zz_AlignerPlugin_logic_extractors_0_maskOh[0];
  assign _zz_AlignerPlugin_logic_extractors_0_maskOh_2 = _zz_AlignerPlugin_logic_extractors_0_maskOh[1];
  assign _zz_AlignerPlugin_logic_extractors_0_maskOh_3 = _zz_AlignerPlugin_logic_extractors_0_maskOh[2];
  always @(*) begin
    _zz_AlignerPlugin_logic_extractors_0_maskOh_4[0] = (_zz_AlignerPlugin_logic_extractors_0_maskOh_1 && (! 1'b0));
    _zz_AlignerPlugin_logic_extractors_0_maskOh_4[1] = (_zz_AlignerPlugin_logic_extractors_0_maskOh_2 && (! _zz_AlignerPlugin_logic_extractors_0_maskOh_1));
    _zz_AlignerPlugin_logic_extractors_0_maskOh_4[2] = (_zz_AlignerPlugin_logic_extractors_0_maskOh_3 && (! ({_zz_AlignerPlugin_logic_extractors_0_maskOh_2,_zz_AlignerPlugin_logic_extractors_0_maskOh_1} != 2'b00)));
    _zz_AlignerPlugin_logic_extractors_0_maskOh_4[3] = (_zz_AlignerPlugin_logic_extractors_0_maskOh[3] && (! ({_zz_AlignerPlugin_logic_extractors_0_maskOh_3,{_zz_AlignerPlugin_logic_extractors_0_maskOh_2,_zz_AlignerPlugin_logic_extractors_0_maskOh_1}} != 3'b000)));
  end

  assign AlignerPlugin_logic_extractors_0_maskOh = _zz_AlignerPlugin_logic_extractors_0_maskOh_4;
  assign _zz_AlignerPlugin_logic_extractors_0_usage = AlignerPlugin_logic_extractors_0_maskOh[0];
  assign _zz_AlignerPlugin_logic_extractors_0_usage_1 = AlignerPlugin_logic_extractors_0_maskOh[1];
  assign _zz_AlignerPlugin_logic_extractors_0_usage_2 = AlignerPlugin_logic_extractors_0_maskOh[2];
  assign _zz_AlignerPlugin_logic_extractors_0_usage_3 = AlignerPlugin_logic_extractors_0_maskOh[3];
  assign AlignerPlugin_logic_extractors_0_usage = (((_zz_AlignerPlugin_logic_extractors_0_usage ? AlignerPlugin_logic_decoders_0_usage : 4'b0000) | (_zz_AlignerPlugin_logic_extractors_0_usage_1 ? AlignerPlugin_logic_decoders_1_usage : 4'b0000)) | ((_zz_AlignerPlugin_logic_extractors_0_usage_2 ? AlignerPlugin_logic_decoders_2_usage : 4'b0000) | (_zz_AlignerPlugin_logic_extractors_0_usage_3 ? AlignerPlugin_logic_decoders_3_usage : 4'b0000)));
  assign AlignerPlugin_logic_extractors_0_usable = _zz_AlignerPlugin_logic_extractors_0_usable[0];
  assign AlignerPlugin_logic_extractors_0_slice0 = (((_zz_AlignerPlugin_logic_extractors_0_usage ? AlignerPlugin_logic_slices_data_0 : 32'h00000000) | (_zz_AlignerPlugin_logic_extractors_0_usage_1 ? AlignerPlugin_logic_slices_data_1 : 32'h00000000)) | ((_zz_AlignerPlugin_logic_extractors_0_usage_2 ? AlignerPlugin_logic_slices_data_2 : 32'h00000000) | (_zz_AlignerPlugin_logic_extractors_0_usage_3 ? AlignerPlugin_logic_slices_data_3 : 32'h00000000)));
  assign AlignerPlugin_logic_extractors_0_valid = ((|AlignerPlugin_logic_slices_carry[3 : 0]) && AlignerPlugin_logic_extractors_0_usable);
  assign FrontendPlugin_aligned_Frontend_INSTRUCTION_ALIGNED_0 = AlignerPlugin_logic_extractors_0_slice0;
  assign FrontendPlugin_aligned_Frontend_MASK_ALIGNED_0 = AlignerPlugin_logic_extractors_0_valid;
  assign AlignerPlugin_logic_extractors_0_sliceLast = FrontendPlugin_aligned_PC_0[2 : 2];
  assign AlignerPlugin_logic_extractors_0_bufferPredictionLast = (AlignerPlugin_logic_buffer_branchSlice == AlignerPlugin_logic_extractors_0_sliceLast);
  assign AlignerPlugin_logic_extractors_0_inputPredictionLast = (AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_SLICE == AlignerPlugin_logic_extractors_0_sliceLast);
  assign AlignerPlugin_logic_extractors_0_lastWord = (|AlignerPlugin_logic_extractors_0_maskOh[3 : 2]);
  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0 = ((AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID && (! _zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1)) && AlignerPlugin_logic_extractors_0_inputPredictionLast);
    end else begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0 = (AlignerPlugin_logic_buffer_branchValid && AlignerPlugin_logic_extractors_0_bufferPredictionLast);
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_0 = AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT;
    end else begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_0 = AlignerPlugin_logic_buffer_branchPcNext;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_BRANCH_HISTORY_0 = AlignerPlugin_setup_s2m_BRANCH_HISTORY;
    end else begin
      FrontendPlugin_aligned_BRANCH_HISTORY_0 = AlignerPlugin_logic_buffer_wordContexts_0;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALID_0 = AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID;
    end else begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALID_0 = AlignerPlugin_logic_buffer_wordContexts_1;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_SLICE_0 = AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_SLICE;
    end else begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_SLICE_0 = AlignerPlugin_logic_buffer_wordContexts_2;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALUE_0 = AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE;
    end else begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALUE_0 = AlignerPlugin_logic_buffer_wordContexts_3;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_GSHARE_COUNTER_0_0 = AlignerPlugin_setup_s2m_GSHARE_COUNTER_0;
    end else begin
      FrontendPlugin_aligned_GSHARE_COUNTER_0_0 = AlignerPlugin_logic_buffer_wordContexts_4_0;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_lastWord) begin
      FrontendPlugin_aligned_GSHARE_COUNTER_0_1 = AlignerPlugin_setup_s2m_GSHARE_COUNTER_1;
    end else begin
      FrontendPlugin_aligned_GSHARE_COUNTER_0_1 = AlignerPlugin_logic_buffer_wordContexts_4_1;
    end
  end

  assign _zz_AlignerPlugin_logic_extractors_0_sliceOffset = AlignerPlugin_logic_extractors_0_maskOh;
  assign _zz_AlignerPlugin_logic_extractors_0_sliceOffset_1 = _zz_AlignerPlugin_logic_extractors_0_sliceOffset[3];
  assign _zz_AlignerPlugin_logic_extractors_0_sliceOffset_2 = (_zz_AlignerPlugin_logic_extractors_0_sliceOffset[1] || _zz_AlignerPlugin_logic_extractors_0_sliceOffset_1);
  assign _zz_AlignerPlugin_logic_extractors_0_sliceOffset_3 = (_zz_AlignerPlugin_logic_extractors_0_sliceOffset[2] || _zz_AlignerPlugin_logic_extractors_0_sliceOffset_1);
  assign AlignerPlugin_logic_extractors_0_sliceOffset = {_zz_AlignerPlugin_logic_extractors_0_sliceOffset_3,_zz_AlignerPlugin_logic_extractors_0_sliceOffset_2};
  assign AlignerPlugin_logic_extractors_0_firstWord = AlignerPlugin_logic_extractors_0_sliceOffset[1];
  assign AlignerPlugin_logic_extractors_0_pcWord = _zz_AlignerPlugin_logic_extractors_0_pcWord;
  assign FrontendPlugin_aligned_PC_0 = {{_zz_FrontendPlugin_aligned_PC_0,AlignerPlugin_logic_extractors_0_sliceOffset[0 : 0]},2'b00};
  always @(*) begin
    if(AlignerPlugin_logic_extractors_0_firstWord) begin
      FrontendPlugin_aligned_FETCH_ID_0 = AlignerPlugin_setup_s2m_FETCH_ID;
    end else begin
      FrontendPlugin_aligned_FETCH_ID_0 = AlignerPlugin_logic_buffer_firstWordContexts_0;
    end
  end

  always @(*) begin
    FrontendPlugin_aligned_Frontend_FETCH_FAULT_0 = 1'b0;
    if(when_AlignerPlugin_l230) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_0 = 1'b1;
    end
    if(when_AlignerPlugin_l235) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_0 = 1'b1;
    end
  end

  always @(*) begin
    FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0 = 1'bx;
    if(when_AlignerPlugin_l230) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0 = AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE;
    end
    if(when_AlignerPlugin_l235) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0 = AlignerPlugin_logic_buffer_fault_page;
    end
  end

  assign when_AlignerPlugin_l230 = ((AlignerPlugin_logic_extractors_0_firstWord || AlignerPlugin_logic_extractors_0_lastWord) && AlignerPlugin_setup_s2m_Fetch_WORD_FAULT);
  assign when_AlignerPlugin_l235 = (((! AlignerPlugin_logic_extractors_0_firstWord) || (! AlignerPlugin_logic_extractors_0_lastWord)) && AlignerPlugin_logic_buffer_fault);
  assign _zz_AlignerPlugin_logic_extractors_1_maskOh = AlignerPlugin_logic_slices_carry_1[3 : 1];
  assign _zz_AlignerPlugin_logic_extractors_1_maskOh_1 = _zz_AlignerPlugin_logic_extractors_1_maskOh[0];
  assign _zz_AlignerPlugin_logic_extractors_1_maskOh_2 = _zz_AlignerPlugin_logic_extractors_1_maskOh[1];
  always @(*) begin
    _zz_AlignerPlugin_logic_extractors_1_maskOh_3[0] = (_zz_AlignerPlugin_logic_extractors_1_maskOh_1 && (! 1'b0));
    _zz_AlignerPlugin_logic_extractors_1_maskOh_3[1] = (_zz_AlignerPlugin_logic_extractors_1_maskOh_2 && (! _zz_AlignerPlugin_logic_extractors_1_maskOh_1));
    _zz_AlignerPlugin_logic_extractors_1_maskOh_3[2] = (_zz_AlignerPlugin_logic_extractors_1_maskOh[2] && (! ({_zz_AlignerPlugin_logic_extractors_1_maskOh_2,_zz_AlignerPlugin_logic_extractors_1_maskOh_1} != 2'b00)));
  end

  assign AlignerPlugin_logic_extractors_1_maskOh = _zz_AlignerPlugin_logic_extractors_1_maskOh_3;
  assign _zz_AlignerPlugin_logic_extractors_1_usage = AlignerPlugin_logic_extractors_1_maskOh[0];
  assign _zz_AlignerPlugin_logic_extractors_1_usage_1 = AlignerPlugin_logic_extractors_1_maskOh[1];
  assign _zz_AlignerPlugin_logic_extractors_1_usage_2 = AlignerPlugin_logic_extractors_1_maskOh[2];
  assign AlignerPlugin_logic_extractors_1_usage = (((_zz_AlignerPlugin_logic_extractors_1_usage ? AlignerPlugin_logic_decoders_1_usage : 4'b0000) | (_zz_AlignerPlugin_logic_extractors_1_usage_1 ? AlignerPlugin_logic_decoders_2_usage : 4'b0000)) | (_zz_AlignerPlugin_logic_extractors_1_usage_2 ? AlignerPlugin_logic_decoders_3_usage : 4'b0000));
  assign AlignerPlugin_logic_extractors_1_usable = _zz_AlignerPlugin_logic_extractors_1_usable[0];
  assign AlignerPlugin_logic_extractors_1_slice0 = (((_zz_AlignerPlugin_logic_extractors_1_usage ? AlignerPlugin_logic_slices_data_1 : 32'h00000000) | (_zz_AlignerPlugin_logic_extractors_1_usage_1 ? AlignerPlugin_logic_slices_data_2 : 32'h00000000)) | (_zz_AlignerPlugin_logic_extractors_1_usage_2 ? AlignerPlugin_logic_slices_data_3 : 32'h00000000));
  always @(*) begin
    AlignerPlugin_logic_extractors_1_valid = ((|AlignerPlugin_logic_slices_carry_1[3 : 1]) && AlignerPlugin_logic_extractors_1_usable);
    if(AlignerPlugin_setup_singleFetch) begin
      AlignerPlugin_logic_extractors_1_valid = 1'b0;
    end
  end

  assign FrontendPlugin_aligned_Frontend_INSTRUCTION_ALIGNED_1 = AlignerPlugin_logic_extractors_1_slice0;
  assign FrontendPlugin_aligned_Frontend_MASK_ALIGNED_1 = AlignerPlugin_logic_extractors_1_valid;
  assign AlignerPlugin_logic_extractors_1_sliceLast = FrontendPlugin_aligned_PC_1[2 : 2];
  assign AlignerPlugin_logic_extractors_1_bufferPredictionLast = (AlignerPlugin_logic_buffer_branchSlice == AlignerPlugin_logic_extractors_1_sliceLast);
  assign AlignerPlugin_logic_extractors_1_inputPredictionLast = (AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_SLICE == AlignerPlugin_logic_extractors_1_sliceLast);
  assign AlignerPlugin_logic_extractors_1_lastWord = (|AlignerPlugin_logic_extractors_1_maskOh[2 : 1]);
  always @(*) begin
    if(AlignerPlugin_logic_extractors_1_lastWord) begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1 = ((AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID && (! _zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1)) && AlignerPlugin_logic_extractors_1_inputPredictionLast);
    end else begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1 = (AlignerPlugin_logic_buffer_branchValid && AlignerPlugin_logic_extractors_1_bufferPredictionLast);
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_1_lastWord) begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_1 = AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT;
    end else begin
      FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_1 = AlignerPlugin_logic_buffer_branchPcNext;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_1_lastWord) begin
      FrontendPlugin_aligned_BRANCH_HISTORY_1 = AlignerPlugin_setup_s2m_BRANCH_HISTORY;
    end else begin
      FrontendPlugin_aligned_BRANCH_HISTORY_1 = AlignerPlugin_logic_buffer_wordContexts_0;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_1_lastWord) begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALID_1 = AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID;
    end else begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALID_1 = AlignerPlugin_logic_buffer_wordContexts_1;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_1_lastWord) begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_SLICE_1 = AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_SLICE;
    end else begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_SLICE_1 = AlignerPlugin_logic_buffer_wordContexts_2;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_1_lastWord) begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALUE_1 = AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE;
    end else begin
      FrontendPlugin_aligned_Prediction_BRANCH_HISTORY_PUSH_VALUE_1 = AlignerPlugin_logic_buffer_wordContexts_3;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_1_lastWord) begin
      FrontendPlugin_aligned_GSHARE_COUNTER_1_0 = AlignerPlugin_setup_s2m_GSHARE_COUNTER_0;
    end else begin
      FrontendPlugin_aligned_GSHARE_COUNTER_1_0 = AlignerPlugin_logic_buffer_wordContexts_4_0;
    end
  end

  always @(*) begin
    if(AlignerPlugin_logic_extractors_1_lastWord) begin
      FrontendPlugin_aligned_GSHARE_COUNTER_1_1 = AlignerPlugin_setup_s2m_GSHARE_COUNTER_1;
    end else begin
      FrontendPlugin_aligned_GSHARE_COUNTER_1_1 = AlignerPlugin_logic_buffer_wordContexts_4_1;
    end
  end

  assign _zz_AlignerPlugin_logic_extractors_1_sliceOffset = ({1'd0,AlignerPlugin_logic_extractors_1_maskOh} <<< 1'd1);
  assign _zz_AlignerPlugin_logic_extractors_1_sliceOffset_1 = _zz_AlignerPlugin_logic_extractors_1_sliceOffset[3];
  assign _zz_AlignerPlugin_logic_extractors_1_sliceOffset_2 = (_zz_AlignerPlugin_logic_extractors_1_sliceOffset[1] || _zz_AlignerPlugin_logic_extractors_1_sliceOffset_1);
  assign _zz_AlignerPlugin_logic_extractors_1_sliceOffset_3 = (_zz_AlignerPlugin_logic_extractors_1_sliceOffset[2] || _zz_AlignerPlugin_logic_extractors_1_sliceOffset_1);
  assign AlignerPlugin_logic_extractors_1_sliceOffset = {_zz_AlignerPlugin_logic_extractors_1_sliceOffset_3,_zz_AlignerPlugin_logic_extractors_1_sliceOffset_2};
  assign AlignerPlugin_logic_extractors_1_firstWord = AlignerPlugin_logic_extractors_1_sliceOffset[1];
  assign AlignerPlugin_logic_extractors_1_pcWord = _zz_AlignerPlugin_logic_extractors_1_pcWord;
  assign FrontendPlugin_aligned_PC_1 = {{_zz_FrontendPlugin_aligned_PC_1,AlignerPlugin_logic_extractors_1_sliceOffset[0 : 0]},2'b00};
  always @(*) begin
    if(AlignerPlugin_logic_extractors_1_firstWord) begin
      FrontendPlugin_aligned_FETCH_ID_1 = AlignerPlugin_setup_s2m_FETCH_ID;
    end else begin
      FrontendPlugin_aligned_FETCH_ID_1 = AlignerPlugin_logic_buffer_firstWordContexts_0;
    end
  end

  always @(*) begin
    FrontendPlugin_aligned_Frontend_FETCH_FAULT_1 = 1'b0;
    if(when_AlignerPlugin_l230_1) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_1 = 1'b1;
    end
    if(when_AlignerPlugin_l235_1) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_1 = 1'b1;
    end
  end

  always @(*) begin
    FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_1 = 1'bx;
    if(when_AlignerPlugin_l230_1) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_1 = AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE;
    end
    if(when_AlignerPlugin_l235_1) begin
      FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_1 = AlignerPlugin_logic_buffer_fault_page;
    end
  end

  assign when_AlignerPlugin_l230_1 = ((AlignerPlugin_logic_extractors_1_firstWord || AlignerPlugin_logic_extractors_1_lastWord) && AlignerPlugin_setup_s2m_Fetch_WORD_FAULT);
  assign when_AlignerPlugin_l235_1 = (((! AlignerPlugin_logic_extractors_1_firstWord) || (! AlignerPlugin_logic_extractors_1_lastWord)) && AlignerPlugin_logic_buffer_fault);
  assign FrontendPlugin_aligned_isFireing = (FrontendPlugin_aligned_valid && FrontendPlugin_aligned_ready);
  assign AlignerPlugin_logic_fireOutput = FrontendPlugin_aligned_isFireing;
  assign AlignerPlugin_logic_fireInput = ((AlignerPlugin_logic_isInputValid && (AlignerPlugin_logic_buffer_mask == 2'b00)) || (AlignerPlugin_logic_fireOutput && (AlignerPlugin_logic_slices_remains_2[1 : 0] == 2'b00)));
  assign AlignerPlugin_logic_postMask = (_zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1 ? 2'b11 : AlignerPlugin_setup_s2m_MASK_BACK);
  assign when_AlignerPlugin_l264 = (AlignerPlugin_setup_s2m_ready || AlignerPlugin_setup_s2m_isFlushed);
  assign _zz_FetchPlugin_stages_1_isFlushingRoot = (_zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1 && (! AlignerPlugin_logic_correctionSent));
  assign AlignerPlugin_setup_sequenceJump_valid = (_zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1 && (! AlignerPlugin_logic_correctionSent));
  assign AlignerPlugin_setup_sequenceJump_payload_pc = AlignerPlugin_setup_s2m_Fetch_FETCH_PC_INC;
  assign FrontendPlugin_aligned_valid = AlignerPlugin_logic_extractors_0_valid;
  assign AlignerPlugin_setup_s2m_haltRequest_AlignerPlugin_l270 = (! AlignerPlugin_logic_fireInput);
  assign FrontendPlugin_decompressed_Frontend_INSTRUCTION_DECOMPRESSED_0 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_0;
  assign FrontendPlugin_decompressed_Frontend_INSTRUCTION_ILLEGAL_0 = 1'b0;
  assign FrontendPlugin_decompressed_Frontend_INSTRUCTION_DECOMPRESSED_1 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_1;
  assign FrontendPlugin_decompressed_Frontend_INSTRUCTION_ILLEGAL_1 = 1'b0;
  assign integer_RfAllocationPlugin_logic_pop_blocked = (! integer_RfAllocationPlugin_logic_allocator_io_pop_ready);
  assign FrontendPlugin_allocated_haltRequest_RfAllocationPlugin_l55 = integer_RfAllocationPlugin_logic_pop_blocked;
  assign when_RfAllocationPlugin_l63 = 1'b1;
  always @(*) begin
    integer_RfAllocationPlugin_logic_allocator_io_pop_mask[0] = ((FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0 && FrontendPlugin_allocated_WRITE_RD_0) && when_RfAllocationPlugin_l63);
    integer_RfAllocationPlugin_logic_allocator_io_pop_mask[1] = ((FrontendPlugin_allocated_Frontend_DISPATCH_MASK_1 && FrontendPlugin_allocated_WRITE_RD_1) && when_RfAllocationPlugin_l63_1);
  end

  always @(*) begin
    FrontendPlugin_allocated_PHYS_RD_0 = 6'bxxxxxx;
    if(when_RfAllocationPlugin_l63) begin
      FrontendPlugin_allocated_PHYS_RD_0 = integer_RfAllocationPlugin_logic_allocator_io_pop_values_0;
    end
  end

  assign when_RfAllocationPlugin_l63_1 = 1'b1;
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RD_1 = 6'bxxxxxx;
    if(when_RfAllocationPlugin_l63_1) begin
      FrontendPlugin_allocated_PHYS_RD_1 = integer_RfAllocationPlugin_logic_allocator_io_pop_values_1;
    end
  end

  assign DispatchPlugin_logic_sparseRob_mask = {FrontendPlugin_serialized_Frontend_DISPATCH_MASK_1,FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0};
  assign DispatchPlugin_logic_sparseRob_remains = (DispatchPlugin_logic_sparseRob_mask & DispatchPlugin_logic_sparseRob_todo);
  assign DispatchPlugin_logic_sparseRob_sparse = ((DispatchPlugin_logic_sparseRob_mask & DispatchPlugin_logic_sparseRob_remains) & {FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_1,FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0});
  assign DispatchPlugin_logic_sparseRob_sparseHit = (|DispatchPlugin_logic_sparseRob_sparse);
  assign DispatchPlugin_logic_sparseRob_sparse_ohFirst_input = DispatchPlugin_logic_sparseRob_sparse;
  assign DispatchPlugin_logic_sparseRob_sparse_ohFirst_masked = (DispatchPlugin_logic_sparseRob_sparse_ohFirst_input & (~ _zz_DispatchPlugin_logic_sparseRob_sparse_ohFirst_masked));
  assign DispatchPlugin_logic_sparseRob_sparseFirst = DispatchPlugin_logic_sparseRob_sparse_ohFirst_masked;
  assign when_DispatchPlugin_l79 = DispatchPlugin_logic_sparseRob_sparse[0];
  always @(*) begin
    if(when_DispatchPlugin_l79) begin
      DispatchPlugin_logic_sparseRob_filter[0] = 1'b1;
    end else begin
      DispatchPlugin_logic_sparseRob_filter[0] = 1'b1;
    end
    if(when_DispatchPlugin_l79_1) begin
      DispatchPlugin_logic_sparseRob_filter[1] = (DispatchPlugin_logic_sparseRob_remains[0 : 0] == 1'b0);
    end else begin
      DispatchPlugin_logic_sparseRob_filter[1] = (DispatchPlugin_logic_sparseRob_sparse[0 : 0] == 1'b0);
    end
  end

  assign when_DispatchPlugin_l79_1 = DispatchPlugin_logic_sparseRob_sparse[1];
  assign DispatchPlugin_logic_sparseRob_masked = (DispatchPlugin_logic_sparseRob_remains & DispatchPlugin_logic_sparseRob_filter);
  assign DispatchPlugin_logic_sparseRob_forkLast = (&(DispatchPlugin_logic_sparseRob_filter | (~ DispatchPlugin_logic_sparseRob_mask)));
  assign FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0_overloaded = (FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0 && DispatchPlugin_logic_sparseRob_masked[0]);
  assign FrontendPlugin_serialized_Frontend_DISPATCH_MASK_1_overloaded = (FrontendPlugin_serialized_Frontend_DISPATCH_MASK_1 && DispatchPlugin_logic_sparseRob_masked[1]);
  assign FrontendPlugin_serialized_forkRequest_DispatchPlugin_l90 = (! DispatchPlugin_logic_sparseRob_forkLast);
  assign when_DispatchPlugin_l94 = (FrontendPlugin_serialized_ready || FrontendPlugin_serialized_isFlushed);
  assign BranchContextPlugin_logic_ptr_occupancy = (BranchContextPlugin_logic_ptr_alloc - BranchContextPlugin_logic_ptr_free);
  assign BranchContextPlugin_logic_alloc_allocNext = BranchContextPlugin_logic_ptr_alloc;
  always @(*) begin
    BranchContextPlugin_logic_alloc_full = 1'b0;
    if(when_BranchContextPlugin_l106) begin
      BranchContextPlugin_logic_alloc_full = 1'b1;
    end
  end

  assign FrontendPlugin_allocated_BRANCH_ID_0 = BranchContextPlugin_logic_alloc_allocNext[3:0];
  assign when_BranchContextPlugin_l93 = ((FrontendPlugin_allocated_valid && FrontendPlugin_allocated_BRANCH_SEL_0) && FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0);
  assign FrontendPlugin_allocated_BRANCH_ID_1 = BranchContextPlugin_logic_alloc_allocNext_1[3:0];
  assign when_BranchContextPlugin_l93_1 = ((FrontendPlugin_allocated_valid && FrontendPlugin_allocated_BRANCH_SEL_1) && FrontendPlugin_allocated_Frontend_DISPATCH_MASK_1);
  assign when_BranchContextPlugin_l106 = (5'h0e < BranchContextPlugin_logic_ptr_occupancy);
  assign FrontendPlugin_allocated_haltRequest_BranchContextPlugin_l107 = BranchContextPlugin_logic_alloc_full;
  always @(*) begin
    DecoderPredictionPlugin_logic_ras_ptr_pushIt = 1'b0;
    if(when_DecoderPredictionPlugin_l212) begin
      DecoderPredictionPlugin_logic_ras_ptr_pushIt = 1'b1;
    end
    if(when_DecoderPredictionPlugin_l212_1) begin
      DecoderPredictionPlugin_logic_ras_ptr_pushIt = 1'b1;
    end
    if(when_DecoderPredictionPlugin_l243) begin
      DecoderPredictionPlugin_logic_ras_ptr_pushIt = 1'b0;
    end
  end

  always @(*) begin
    DecoderPredictionPlugin_logic_ras_ptr_popIt = 1'b0;
    if(when_DecoderPredictionPlugin_l219) begin
      DecoderPredictionPlugin_logic_ras_ptr_popIt = 1'b1;
    end
    if(when_DecoderPredictionPlugin_l219_1) begin
      DecoderPredictionPlugin_logic_ras_ptr_popIt = 1'b1;
    end
    if(when_DecoderPredictionPlugin_l244) begin
      DecoderPredictionPlugin_logic_ras_ptr_popIt = 1'b0;
    end
  end

  assign DecoderPredictionPlugin_logic_ras_read = _zz_DecoderPredictionPlugin_logic_ras_mem_stack_port0;
  assign DecoderPredictionPlugin_logic_ras_write_valid = DecoderPredictionPlugin_logic_ras_ptr_pushIt;
  assign DecoderPredictionPlugin_logic_ras_write_payload_address = DecoderPredictionPlugin_logic_ras_ptr_push;
  always @(*) begin
    DecoderPredictionPlugin_logic_ras_write_payload_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_DecoderPredictionPlugin_l212) begin
      if(when_DecoderPredictionPlugin_l213) begin
        DecoderPredictionPlugin_logic_ras_write_payload_data = FrontendPlugin_serialized_PC_INC_0;
      end
    end
    if(when_DecoderPredictionPlugin_l212_1) begin
      if(when_DecoderPredictionPlugin_l213_1) begin
        DecoderPredictionPlugin_logic_ras_write_payload_data = FrontendPlugin_serialized_PC_INC_1;
      end
    end
  end

  assign BtbPlugin_logic_onLearn_hash = BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[18 : 3];
  assign BtbPlugin_logic_onLearn_port_valid = BranchContextPlugin_setup_learnValid;
  assign BtbPlugin_logic_onLearn_port_payload_address = _zz_BtbPlugin_logic_onLearn_port_payload_address[8:0];
  assign BtbPlugin_logic_onLearn_port_payload_data_hash = BtbPlugin_logic_onLearn_hash;
  assign BtbPlugin_logic_onLearn_port_payload_data_slice = _zz_BtbPlugin_logic_onLearn_port_payload_data_slice[0:0];
  assign BtbPlugin_logic_onLearn_port_payload_data_pcTarget = BranchContextPlugin_learn_BRANCH_FINAL_pcTarget;
  assign BtbPlugin_logic_onLearn_port_payload_data_isBranch = BranchContextPlugin_free_learn_Prediction_IS_BRANCH;
  assign BtbPlugin_logic_readCmd_entryAddress = _zz_BtbPlugin_logic_readCmd_entryAddress[8:0];
  assign _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash = _zz_BtbPlugin_logic_mem_port1;
  assign FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash = _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash[15 : 0];
  assign FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_slice = _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash[16 : 16];
  assign FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_pcTarget = _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash[48 : 17];
  assign FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_isBranch = _zz_FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash[49];
  assign BtbPlugin_logic_hitCalc_postPcPrediction = (FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_slice < FetchPlugin_stages_1_Fetch_FETCH_PC[2 : 2]);
  assign FetchPlugin_stages_1_BtbPlugin_logic_HIT = ((FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_hash == FetchPlugin_stages_1_Fetch_FETCH_PC[18 : 3]) && (! BtbPlugin_logic_hitCalc_postPcPrediction));
  assign BtbPlugin_logic_applyIt_prediction = _zz_BtbPlugin_logic_applyIt_prediction;
  assign BtbPlugin_logic_applyIt_needIt = ((FetchPlugin_stages_1_valid && FetchPlugin_stages_1_BtbPlugin_logic_HIT) && (! (FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_isBranch && (! BtbPlugin_logic_applyIt_prediction))));
  assign when_BtbPlugin_l109 = (FetchPlugin_stages_1_ready || FetchPlugin_stages_1_isFlushed);
  assign BtbPlugin_logic_applyIt_doIt = (BtbPlugin_logic_applyIt_needIt && (! BtbPlugin_logic_applyIt_correctionSent));
  assign BtbPlugin_setup_btbJump_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_setup_btbJump_payload_pc = FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_pcTarget;
  assign FetchPlugin_stages_1_Prediction_WORD_BRANCH_VALID = BtbPlugin_logic_applyIt_needIt;
  assign FetchPlugin_stages_1_Prediction_WORD_BRANCH_SLICE = FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_slice;
  assign FetchPlugin_stages_1_Prediction_WORD_BRANCH_PC_NEXT = FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_pcTarget;
  assign BtbPlugin_setup_historyPush_flush = (((FetchPlugin_stages_1_valid && FetchPlugin_stages_1_BtbPlugin_logic_HIT) && FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_isBranch) && (! BtbPlugin_logic_applyIt_correctionSent));
  assign BtbPlugin_setup_historyPush_mask[0] = BtbPlugin_setup_historyPush_flush;
  assign BtbPlugin_setup_historyPush_taken[0] = BtbPlugin_logic_applyIt_prediction;
  assign FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALID = BtbPlugin_setup_historyPush_flush;
  assign FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_SLICE = FetchPlugin_stages_1_BtbPlugin_logic_ENTRY_slice;
  assign FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALUE = BtbPlugin_logic_applyIt_prediction;
  assign _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH = FetchPlugin_stages_0_Fetch_FETCH_PC[15 : 3];
  assign FetchPlugin_stages_0_GSharePlugin_logic_HASH = ({_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[0],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[1],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[2],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[3],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[4],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH[5],{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_1,{_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_2,_zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_3}}}}}}}} ^ _zz_FetchPlugin_stages_0_GSharePlugin_logic_HASH_4);
  assign FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_valid = GSharePlugin_logic_mem_write_valid;
  assign FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_address = GSharePlugin_logic_mem_write_payload_address;
  assign FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_data_0 = GSharePlugin_logic_mem_write_payload_data_0;
  assign FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_data_1 = GSharePlugin_logic_mem_write_payload_data_1;
  assign _zz_FetchPlugin_stages_1_GSHARE_COUNTER_0 = _zz_FetchPlugin_stages_1_GSHARE_COUNTER_0_1;
  always @(*) begin
    FetchPlugin_stages_1_GSHARE_COUNTER_0 = _zz_FetchPlugin_stages_1_GSHARE_COUNTER_0[1 : 0];
    if(when_GSharePlugin_l98) begin
      FetchPlugin_stages_1_GSHARE_COUNTER_0 = FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_data_0;
    end
  end

  always @(*) begin
    FetchPlugin_stages_1_GSHARE_COUNTER_1 = _zz_FetchPlugin_stages_1_GSHARE_COUNTER_0[3 : 2];
    if(when_GSharePlugin_l98) begin
      FetchPlugin_stages_1_GSHARE_COUNTER_1 = FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_data_1;
    end
  end

  assign when_GSharePlugin_l98 = (FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_valid && (FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_address == FetchPlugin_stages_1_GSharePlugin_logic_HASH));
  assign FrontendPlugin_decompressed_Prediction_CONDITIONAL_TAKE_IT_0 = {FrontendPlugin_decompressed_GSHARE_COUNTER_0_1[1],FrontendPlugin_decompressed_GSHARE_COUNTER_0_0[1]};
  assign FrontendPlugin_decompressed_Prediction_CONDITIONAL_TAKE_IT_1 = {FrontendPlugin_decompressed_GSHARE_COUNTER_1_1[1],FrontendPlugin_decompressed_GSHARE_COUNTER_1_0[1]};
  assign _zz_GSharePlugin_logic_onLearn_hash = BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[15 : 3];
  assign GSharePlugin_logic_onLearn_hash = ({_zz_GSharePlugin_logic_onLearn_hash[0],{_zz_GSharePlugin_logic_onLearn_hash[1],{_zz_GSharePlugin_logic_onLearn_hash[2],{_zz_GSharePlugin_logic_onLearn_hash[3],{_zz_GSharePlugin_logic_onLearn_hash[4],{_zz_GSharePlugin_logic_onLearn_hash[5],{_zz_GSharePlugin_logic_onLearn_hash_1,{_zz_GSharePlugin_logic_onLearn_hash_2,_zz_GSharePlugin_logic_onLearn_hash_3}}}}}}}} ^ _zz_GSharePlugin_logic_onLearn_hash_4);
  assign GSharePlugin_logic_onLearn_incrValue = (BranchContextPlugin_learn_BRANCH_FINAL_taken ? 2'b01 : 2'b11);
  always @(*) begin
    GSharePlugin_logic_onLearn_overflow = 1'b0;
    if(when_GSharePlugin_l123) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
    if(when_GSharePlugin_l123_1) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
  end

  assign GSharePlugin_logic_onLearn_updated_0 = (BranchContextPlugin_free_learn_GSHARE_COUNTER_0 + ((BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[2 : 2] == 1'b0) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l123 = (((BranchContextPlugin_learn_BRANCH_FINAL_taken && BranchContextPlugin_free_learn_GSHARE_COUNTER_0[1]) && (! GSharePlugin_logic_onLearn_updated_0[1])) || (((! BranchContextPlugin_learn_BRANCH_FINAL_taken) && (! BranchContextPlugin_free_learn_GSHARE_COUNTER_0[1])) && GSharePlugin_logic_onLearn_updated_0[1]));
  assign GSharePlugin_logic_onLearn_updated_1 = (BranchContextPlugin_free_learn_GSHARE_COUNTER_1 + ((BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[2 : 2] == 1'b1) ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l123_1 = (((BranchContextPlugin_learn_BRANCH_FINAL_taken && BranchContextPlugin_free_learn_GSHARE_COUNTER_1[1]) && (! GSharePlugin_logic_onLearn_updated_1[1])) || (((! BranchContextPlugin_learn_BRANCH_FINAL_taken) && (! BranchContextPlugin_free_learn_GSHARE_COUNTER_1[1])) && GSharePlugin_logic_onLearn_updated_1[1]));
  assign GSharePlugin_logic_mem_write_valid = ((BranchContextPlugin_setup_learnValid && BranchContextPlugin_free_learn_Prediction_IS_BRANCH) && (! GSharePlugin_logic_onLearn_overflow));
  assign GSharePlugin_logic_mem_write_payload_address = GSharePlugin_logic_onLearn_hash;
  assign GSharePlugin_logic_mem_write_payload_data_0 = GSharePlugin_logic_onLearn_updated_0;
  assign GSharePlugin_logic_mem_write_payload_data_1 = GSharePlugin_logic_onLearn_updated_1;
  assign DataCachePlugin_setup_writebackBusy = DataCachePlugin_logic_cache_io_writebackBusy;
  assign DataCachePlugin_setup_refillEvent = toplevel_DataCachePlugin_logic_cache_io_refillEvent_regNext;
  assign DataCachePlugin_setup_writebackEvent = toplevel_DataCachePlugin_logic_cache_io_writebackEvent_regNext;
  assign DataCachePlugin_setup_refillCompletions = DataCachePlugin_logic_cache_io_refillCompletions;
  assign DataCachePlugin_logic_load_hits = {Lsu2Plugin_setup_cacheLoad_cmd_valid,MmuPlugin_setup_cacheLoad_cmd_valid};
  assign DataCachePlugin_logic_load_hit = (|DataCachePlugin_logic_load_hits);
  assign _zz_DataCachePlugin_logic_load_hits_bools_0 = DataCachePlugin_logic_load_hits;
  assign DataCachePlugin_logic_load_hits_bools_0 = _zz_DataCachePlugin_logic_load_hits_bools_0[0];
  assign DataCachePlugin_logic_load_hits_bools_1 = _zz_DataCachePlugin_logic_load_hits_bools_0[1];
  always @(*) begin
    _zz_DataCachePlugin_logic_load_oh[0] = (DataCachePlugin_logic_load_hits_bools_0 && (! 1'b0));
    _zz_DataCachePlugin_logic_load_oh[1] = (DataCachePlugin_logic_load_hits_bools_1 && (! DataCachePlugin_logic_load_hits_bools_0));
  end

  assign DataCachePlugin_logic_load_oh = _zz_DataCachePlugin_logic_load_oh;
  assign _zz_DataCachePlugin_logic_load_ohHistory_0 = DataCachePlugin_logic_load_oh;
  assign DataCachePlugin_logic_load_ohHistory_0 = _zz_DataCachePlugin_logic_load_ohHistory_0;
  assign DataCachePlugin_logic_load_ohHistory_1 = _zz_DataCachePlugin_logic_load_ohHistory_1;
  assign DataCachePlugin_logic_load_ohHistory_2 = _zz_DataCachePlugin_logic_load_ohHistory_2;
  assign _zz_MmuPlugin_setup_cacheLoad_cmd_ready = DataCachePlugin_logic_load_oh[0];
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_virtual = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_virtual : Lsu2Plugin_setup_cacheLoad_cmd_payload_virtual);
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_size = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_size : Lsu2Plugin_setup_cacheLoad_cmd_payload_size);
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_redoOnDataHazard = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_redoOnDataHazard : Lsu2Plugin_setup_cacheLoad_cmd_payload_redoOnDataHazard);
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_unlocked = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_unlocked : Lsu2Plugin_setup_cacheLoad_cmd_payload_unlocked);
  assign DataCachePlugin_logic_cache_io_load_cmd_payload_unique = (_zz_MmuPlugin_setup_cacheLoad_cmd_ready ? MmuPlugin_setup_cacheLoad_cmd_payload_unique : Lsu2Plugin_setup_cacheLoad_cmd_payload_unique);
  assign MmuPlugin_setup_cacheLoad_cmd_ready = _zz_MmuPlugin_setup_cacheLoad_cmd_ready;
  assign Lsu2Plugin_setup_cacheLoad_cmd_ready = DataCachePlugin_logic_load_oh[1];
  assign DataCachePlugin_logic_cache_io_load_cancels = (MmuPlugin_setup_cacheLoad_cancels | Lsu2Plugin_setup_cacheLoad_cancels);
  assign _zz_io_load_translated_physical = DataCachePlugin_logic_load_ohHistory_1[0];
  assign DataCachePlugin_logic_cache_io_load_translated_physical = (_zz_io_load_translated_physical ? MmuPlugin_setup_cacheLoad_translated_physical : Lsu2Plugin_setup_cacheLoad_translated_physical);
  assign DataCachePlugin_logic_cache_io_load_translated_abord = (_zz_io_load_translated_physical ? MmuPlugin_setup_cacheLoad_translated_abord : Lsu2Plugin_setup_cacheLoad_translated_abord);
  assign MmuPlugin_setup_cacheLoad_rsp_valid = (DataCachePlugin_logic_cache_io_load_rsp_valid && DataCachePlugin_logic_load_ohHistory_2[0]);
  assign MmuPlugin_setup_cacheLoad_rsp_payload_data = DataCachePlugin_logic_cache_io_load_rsp_payload_data;
  assign MmuPlugin_setup_cacheLoad_rsp_payload_fault = DataCachePlugin_logic_cache_io_load_rsp_payload_fault;
  assign MmuPlugin_setup_cacheLoad_rsp_payload_redo = DataCachePlugin_logic_cache_io_load_rsp_payload_redo;
  assign MmuPlugin_setup_cacheLoad_rsp_payload_refillSlot = DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlot;
  assign MmuPlugin_setup_cacheLoad_rsp_payload_refillSlotAny = DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlotAny;
  assign Lsu2Plugin_setup_cacheLoad_rsp_valid = (DataCachePlugin_logic_cache_io_load_rsp_valid && DataCachePlugin_logic_load_ohHistory_2[1]);
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_data = DataCachePlugin_logic_cache_io_load_rsp_payload_data;
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_fault = DataCachePlugin_logic_cache_io_load_rsp_payload_fault;
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_redo = DataCachePlugin_logic_cache_io_load_rsp_payload_redo;
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlot = DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlot;
  assign Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlotAny = DataCachePlugin_logic_cache_io_load_rsp_payload_refillSlotAny;
  assign Lsu2Plugin_setup_cacheStore_cmd_ready = DataCachePlugin_logic_cache_io_store_cmd_ready;
  assign Lsu2Plugin_setup_cacheStore_rsp_valid = DataCachePlugin_logic_cache_io_store_rsp_valid;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_fault = DataCachePlugin_logic_cache_io_store_rsp_payload_fault;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_redo = DataCachePlugin_logic_cache_io_store_rsp_payload_redo;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlot = DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlot;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlotAny = DataCachePlugin_logic_cache_io_store_rsp_payload_refillSlotAny;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_generationKo = DataCachePlugin_logic_cache_io_store_rsp_payload_generationKo;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_flush = DataCachePlugin_logic_cache_io_store_rsp_payload_flush;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_prefetch = DataCachePlugin_logic_cache_io_store_rsp_payload_prefetch;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_address = DataCachePlugin_logic_cache_io_store_rsp_payload_address;
  assign Lsu2Plugin_setup_cacheStore_rsp_payload_io = DataCachePlugin_logic_cache_io_store_rsp_payload_io;
  assign DataCachePlugin_mem_read_cmd_valid = DataCachePlugin_logic_cache_io_mem_read_cmd_valid;
  assign DataCachePlugin_mem_read_cmd_payload_id = DataCachePlugin_logic_cache_io_mem_read_cmd_payload_id;
  assign DataCachePlugin_mem_read_cmd_payload_address = DataCachePlugin_logic_cache_io_mem_read_cmd_payload_address;
  assign DataCachePlugin_mem_read_rsp_ready = DataCachePlugin_logic_cache_io_mem_read_rsp_ready;
  assign DataCachePlugin_mem_write_cmd_valid = DataCachePlugin_logic_cache_io_mem_write_cmd_valid;
  assign DataCachePlugin_mem_write_cmd_payload_last = DataCachePlugin_logic_cache_io_mem_write_cmd_payload_last;
  assign DataCachePlugin_mem_write_cmd_payload_fragment_address = DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_address;
  assign DataCachePlugin_mem_write_cmd_payload_fragment_data = DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_data;
  assign DataCachePlugin_mem_write_cmd_payload_fragment_id = DataCachePlugin_logic_cache_io_mem_write_cmd_payload_fragment_id;
  assign CommitPlugin_logic_ptr_commitRow = (CommitPlugin_logic_ptr_commit >>> 1'd1);
  always @(*) begin
    CommitPlugin_logic_ptr_commitNext = CommitPlugin_logic_ptr_commit;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_logic_commit_lineCommited) begin
        CommitPlugin_logic_ptr_commitNext = (CommitPlugin_logic_ptr_commit + 7'h02);
      end
      if(CommitPlugin_logic_commit_rescheduleHit) begin
        CommitPlugin_logic_ptr_commitNext = CommitPlugin_logic_ptr_allocNext;
      end
    end
  end

  assign CommitPlugin_logic_ptr_full = ((CommitPlugin_logic_ptr_alloc ^ CommitPlugin_logic_ptr_free) == 7'h40);
  assign CommitPlugin_logic_ptr_canFree = (CommitPlugin_logic_ptr_free != CommitPlugin_logic_ptr_commit);
  assign CommitPlugin_setup_robLineMask_line = CommitPlugin_logic_ptr_commitNext[5:0];
  assign FrontendPlugin_allocated_ROB_ID = CommitPlugin_logic_ptr_alloc[5:0];
  assign FrontendPlugin_allocated_ROB_MSB_0 = CommitPlugin_logic_ptr_alloc[6];
  assign FrontendPlugin_allocated_ROB_MSB_1 = CommitPlugin_logic_ptr_alloc[6];
  assign FrontendPlugin_allocated_haltRequest_CommitPlugin_l95 = CommitPlugin_logic_ptr_full;
  assign CommitPlugin_logic_ptr_allocNext = (CommitPlugin_logic_ptr_alloc + _zz_CommitPlugin_logic_ptr_allocNext);
  assign CommitPlugin_setup_isRobEmpty = CommitPlugin_logic_ptr_empty;
  assign CommitPlugin_logic_reschedule_commit_row = CommitPlugin_logic_reschedule_robId[5 : 1];
  assign CommitPlugin_logic_reschedule_commit_col = CommitPlugin_logic_reschedule_robId[0 : 0];
  assign CommitPlugin_logic_reschedule_commit_rowHit = (CommitPlugin_logic_reschedule_valid && (CommitPlugin_logic_reschedule_commit_row == _zz_CommitPlugin_logic_reschedule_commit_rowHit));
  assign CommitPlugin_logic_reschedule_age = (CommitPlugin_logic_reschedule_robId - _zz_CommitPlugin_logic_reschedule_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_0_age = (Lsu2Plugin_setup_sharedTrap_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_0_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_1_age = (Lsu2Plugin_setup_specialTrap_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_1_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_2_age = (ALU0_BranchPlugin_setup_reschedule_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_2_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_3_age = (EnvCallPlugin_setup_reschedule_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_3_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_4_age = (EU0_CsrAccessPlugin_setup_trap_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_4_age);
  assign CommitPlugin_logic_reschedule_portsLogic_perPort_5_age = (ALU1_BranchPlugin_setup_reschedule_payload_robId - _zz_CommitPlugin_logic_reschedule_portsLogic_perPort_5_age);
  always @(*) begin
    CommitPlugin_logic_reschedule_portsLogic_hits[0] = (Lsu2Plugin_setup_sharedTrap_valid && ((((((_zz_CommitPlugin_logic_reschedule_portsLogic_hits || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_1) && (_zz_CommitPlugin_logic_reschedule_portsLogic_hits_2 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_3)) && ((! ALU0_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_2_age))) && ((! EnvCallPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_3_age))) && ((! EU0_CsrAccessPlugin_setup_trap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_4_age))) && ((! ALU1_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_0_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_5_age))));
    CommitPlugin_logic_reschedule_portsLogic_hits[1] = (Lsu2Plugin_setup_specialTrap_valid && ((((((_zz_CommitPlugin_logic_reschedule_portsLogic_hits_4 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_5) && (_zz_CommitPlugin_logic_reschedule_portsLogic_hits_6 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_7)) && ((! ALU0_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_2_age))) && ((! EnvCallPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_3_age))) && ((! EU0_CsrAccessPlugin_setup_trap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_4_age))) && ((! ALU1_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_1_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_5_age))));
    CommitPlugin_logic_reschedule_portsLogic_hits[2] = (ALU0_BranchPlugin_setup_reschedule_valid && (((((((! CommitPlugin_logic_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age < CommitPlugin_logic_reschedule_age)) && ((! Lsu2Plugin_setup_sharedTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age < CommitPlugin_logic_reschedule_portsLogic_perPort_0_age))) && ((! Lsu2Plugin_setup_specialTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age < CommitPlugin_logic_reschedule_portsLogic_perPort_1_age))) && ((! EnvCallPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_3_age))) && ((! EU0_CsrAccessPlugin_setup_trap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_4_age))) && ((! ALU1_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_2_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_5_age))));
    CommitPlugin_logic_reschedule_portsLogic_hits[3] = (EnvCallPlugin_setup_reschedule_valid && ((((((_zz_CommitPlugin_logic_reschedule_portsLogic_hits_8 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_9) && (_zz_CommitPlugin_logic_reschedule_portsLogic_hits_10 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_11)) && ((! Lsu2Plugin_setup_specialTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age < CommitPlugin_logic_reschedule_portsLogic_perPort_1_age))) && ((! ALU0_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age < CommitPlugin_logic_reschedule_portsLogic_perPort_2_age))) && ((! EU0_CsrAccessPlugin_setup_trap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_4_age))) && ((! ALU1_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_3_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_5_age))));
    CommitPlugin_logic_reschedule_portsLogic_hits[4] = (EU0_CsrAccessPlugin_setup_trap_valid && ((((((_zz_CommitPlugin_logic_reschedule_portsLogic_hits_12 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_13) && (_zz_CommitPlugin_logic_reschedule_portsLogic_hits_14 || _zz_CommitPlugin_logic_reschedule_portsLogic_hits_15)) && ((! Lsu2Plugin_setup_specialTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_portsLogic_perPort_1_age))) && ((! ALU0_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_portsLogic_perPort_2_age))) && ((! EnvCallPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age < CommitPlugin_logic_reschedule_portsLogic_perPort_3_age))) && ((! ALU1_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_4_age <= CommitPlugin_logic_reschedule_portsLogic_perPort_5_age))));
    CommitPlugin_logic_reschedule_portsLogic_hits[5] = (ALU1_BranchPlugin_setup_reschedule_valid && (((((((! CommitPlugin_logic_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_5_age < CommitPlugin_logic_reschedule_age)) && ((! Lsu2Plugin_setup_sharedTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_5_age < CommitPlugin_logic_reschedule_portsLogic_perPort_0_age))) && ((! Lsu2Plugin_setup_specialTrap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_5_age < CommitPlugin_logic_reschedule_portsLogic_perPort_1_age))) && ((! ALU0_BranchPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_5_age < CommitPlugin_logic_reschedule_portsLogic_perPort_2_age))) && ((! EnvCallPlugin_setup_reschedule_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_5_age < CommitPlugin_logic_reschedule_portsLogic_perPort_3_age))) && ((! EU0_CsrAccessPlugin_setup_trap_valid) || (CommitPlugin_logic_reschedule_portsLogic_perPort_5_age < CommitPlugin_logic_reschedule_portsLogic_perPort_4_age))));
  end

  assign when_CommitPlugin_l131 = (|CommitPlugin_logic_reschedule_portsLogic_hits);
  assign _zz_CommitPlugin_logic_reschedule_trap = CommitPlugin_logic_reschedule_portsLogic_hits[0];
  assign _zz_CommitPlugin_logic_reschedule_trap_1 = CommitPlugin_logic_reschedule_portsLogic_hits[1];
  assign _zz_CommitPlugin_logic_reschedule_trap_2 = CommitPlugin_logic_reschedule_portsLogic_hits[2];
  assign _zz_CommitPlugin_logic_reschedule_trap_3 = CommitPlugin_logic_reschedule_portsLogic_hits[3];
  assign _zz_CommitPlugin_logic_reschedule_trap_4 = CommitPlugin_logic_reschedule_portsLogic_hits[4];
  assign _zz_CommitPlugin_logic_reschedule_trap_5 = CommitPlugin_logic_reschedule_portsLogic_hits[5];
  assign CommitPlugin_setup_jump_valid = (CommitPlugin_logic_reschedule_fresh && (! CommitPlugin_logic_reschedule_trap));
  assign CommitPlugin_setup_jump_payload_pc = CommitPlugin_logic_reschedule_pcTarget;
  assign CommitPlugin_logic_reschedule_reschedulePort_valid = CommitPlugin_logic_reschedule_fresh;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_robId = CommitPlugin_logic_reschedule_robId;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_trap = CommitPlugin_logic_reschedule_trap;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_cause = CommitPlugin_logic_reschedule_cause;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_tval = CommitPlugin_logic_reschedule_tval;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_reason = CommitPlugin_logic_reschedule_reason;
  assign CommitPlugin_logic_reschedule_reschedulePort_payload_skipCommit = CommitPlugin_logic_reschedule_skipCommit;
  always @(*) begin
    CommitPlugin_logic_commit_rescheduleHit = 1'b0;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_commit_slot_0_enable) begin
        if(CommitPlugin_logic_commit_continue) begin
          if(when_CommitPlugin_l207) begin
            CommitPlugin_logic_commit_rescheduleHit = 1'b1;
          end
        end
      end
      if(CommitPlugin_commit_slot_1_enable) begin
        if(CommitPlugin_logic_commit_continue_1) begin
          if(when_CommitPlugin_l207_1) begin
            CommitPlugin_logic_commit_rescheduleHit = 1'b1;
          end
        end
      end
    end
  end

  assign CommitPlugin_logic_commit_active = {_zz_CommitPlugin_logic_commit_active_2[1],_zz_CommitPlugin_logic_commit_active_2[0]};
  always @(*) begin
    CommitPlugin_logic_commit_maskComb = CommitPlugin_logic_commit_mask;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_commit_slot_0_enable) begin
        if(CommitPlugin_logic_commit_continue) begin
          if(when_CommitPlugin_l203) begin
            CommitPlugin_logic_commit_maskComb[0] = 1'b0;
          end
        end
      end
      if(CommitPlugin_commit_slot_1_enable) begin
        if(CommitPlugin_logic_commit_continue_1) begin
          if(when_CommitPlugin_l203_1) begin
            CommitPlugin_logic_commit_maskComb[1] = 1'b0;
          end
        end
      end
    end
  end

  assign CommitPlugin_logic_commit_lineCommited = ((CommitPlugin_logic_commit_maskComb & CommitPlugin_logic_commit_active) == 2'b00);
  always @(*) begin
    CommitPlugin_logic_commit_event_mask = 2'b00;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_commit_slot_0_enable) begin
        if(CommitPlugin_logic_commit_continue) begin
          if(when_CommitPlugin_l203) begin
            CommitPlugin_logic_commit_event_mask[0] = 1'b1;
          end
        end
      end
      if(CommitPlugin_commit_slot_1_enable) begin
        if(CommitPlugin_logic_commit_continue_1) begin
          if(when_CommitPlugin_l203_1) begin
            CommitPlugin_logic_commit_event_mask[1] = 1'b1;
          end
        end
      end
    end
  end

  assign CommitPlugin_logic_commit_event_robId = CommitPlugin_logic_ptr_commit[5:0];
  always @(*) begin
    CommitPlugin_logic_commit_lineEvent_valid = 1'b0;
    if(when_CommitPlugin_l194) begin
      if(when_CommitPlugin_l217) begin
        CommitPlugin_logic_commit_lineEvent_valid = 1'b1;
      end
    end
  end

  assign CommitPlugin_logic_commit_lineEvent_payload_mask = (CommitPlugin_logic_commit_active ^ CommitPlugin_logic_commit_maskComb);
  assign CommitPlugin_logic_commit_lineEvent_payload_robId = CommitPlugin_logic_ptr_commit[5:0];
  assign CommitPlugin_logic_commit_reschedulePort_valid = CommitPlugin_logic_commit_rescheduleHit;
  assign CommitPlugin_logic_commit_reschedulePort_payload_robId = CommitPlugin_logic_reschedule_robId;
  assign CommitPlugin_logic_commit_reschedulePort_payload_robIdNext = CommitPlugin_logic_ptr_allocNext[5:0];
  assign CommitPlugin_logic_commit_reschedulePort_payload_trap = CommitPlugin_logic_reschedule_trap;
  assign CommitPlugin_logic_commit_reschedulePort_payload_cause = CommitPlugin_logic_reschedule_cause;
  assign CommitPlugin_logic_commit_reschedulePort_payload_tval = CommitPlugin_logic_reschedule_tval;
  assign CommitPlugin_logic_commit_reschedulePort_payload_reason = CommitPlugin_logic_reschedule_reason;
  assign CommitPlugin_logic_commit_reschedulePort_payload_skipCommit = CommitPlugin_logic_reschedule_skipCommit;
  always @(*) begin
    CommitPlugin_logic_commit_headNext = CommitPlugin_logic_commit_head;
    if(when_CommitPlugin_l194) begin
      if(CommitPlugin_logic_commit_rescheduleHit) begin
        CommitPlugin_logic_commit_headNext = CommitPlugin_logic_ptr_allocNext[5:0];
      end
    end
  end

  assign _zz_CommitPlugin_logic_commit_head = (CommitPlugin_logic_commit_active & CommitPlugin_logic_commit_mask);
  assign _zz_CommitPlugin_logic_commit_head_1 = _zz__zz_CommitPlugin_logic_commit_head_1[1];
  assign CommitPlugin_logic_commit_head = _zz_CommitPlugin_logic_commit_head_2[5:0];
  assign CommitPlugin_logic_commit_continue = 1'b1;
  assign when_CommitPlugin_l194 = (! CommitPlugin_logic_ptr_empty);
  assign CommitPlugin_commit_slot_0_enable = (CommitPlugin_logic_commit_mask[0] && CommitPlugin_logic_commit_active[0]);
  assign CommitPlugin_commit_slot_0_readyForCommit = CommitPlugin_logic_ptr_robLineMaskRsp[0];
  assign CommitPlugin_commit_slot_0_rescheduleHitSlot = (CommitPlugin_logic_reschedule_commit_rowHit && (CommitPlugin_logic_reschedule_commit_col == 1'b0));
  assign when_CommitPlugin_l203 = (CommitPlugin_commit_slot_0_readyForCommit && (! (CommitPlugin_commit_slot_0_rescheduleHitSlot && CommitPlugin_logic_reschedule_skipCommit)));
  assign when_CommitPlugin_l207 = (CommitPlugin_commit_slot_0_rescheduleHitSlot && (CommitPlugin_logic_reschedule_skipCommit || CommitPlugin_commit_slot_0_readyForCommit));
  assign when_CommitPlugin_l211 = ((! CommitPlugin_commit_slot_0_readyForCommit) || CommitPlugin_commit_slot_0_rescheduleHitSlot);
  assign CommitPlugin_commit_slot_1_enable = (CommitPlugin_logic_commit_mask[1] && CommitPlugin_logic_commit_active[1]);
  assign CommitPlugin_commit_slot_1_readyForCommit = CommitPlugin_logic_ptr_robLineMaskRsp[1];
  assign CommitPlugin_commit_slot_1_rescheduleHitSlot = (CommitPlugin_logic_reschedule_commit_rowHit && (CommitPlugin_logic_reschedule_commit_col == 1'b1));
  assign when_CommitPlugin_l203_1 = (CommitPlugin_commit_slot_1_readyForCommit && (! (CommitPlugin_commit_slot_1_rescheduleHitSlot && CommitPlugin_logic_reschedule_skipCommit)));
  assign when_CommitPlugin_l207_1 = (CommitPlugin_commit_slot_1_rescheduleHitSlot && (CommitPlugin_logic_reschedule_skipCommit || CommitPlugin_commit_slot_1_readyForCommit));
  assign when_CommitPlugin_l211_1 = ((! CommitPlugin_commit_slot_1_readyForCommit) || CommitPlugin_commit_slot_1_rescheduleHitSlot);
  assign when_CommitPlugin_l217 = (CommitPlugin_logic_commit_lineCommited || CommitPlugin_logic_commit_rescheduleHit);
  assign CommitPlugin_logic_free_lineEventStream_valid = CommitPlugin_logic_commit_lineEvent_valid;
  assign CommitPlugin_logic_free_lineEventStream_payload_robId = CommitPlugin_logic_commit_lineEvent_payload_robId;
  assign CommitPlugin_logic_free_lineEventStream_payload_mask = CommitPlugin_logic_commit_lineEvent_payload_mask;
  assign CommitPlugin_logic_free_lineEventStream_ready = CommitPlugin_logic_free_lineEventStream_fifo_io_push_ready;
  assign CommitPlugin_logic_free_robHit = (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_robId == _zz_CommitPlugin_logic_free_robHit);
  assign CommitPlugin_logic_free_hit = (CommitPlugin_logic_free_lineEventStream_fifo_io_pop_valid && CommitPlugin_logic_free_robHit);
  assign CommitPlugin_logic_free_lineEventStream_fifo_io_pop_ready = (CommitPlugin_logic_free_robHit && CommitPlugin_logic_ptr_canFree);
  assign CommitPlugin_logic_free_port_valid = CommitPlugin_logic_ptr_canFree;
  assign CommitPlugin_logic_free_port_payload_robId = CommitPlugin_logic_ptr_free[5:0];
  assign CommitPlugin_logic_free_port_payload_commited = (CommitPlugin_logic_free_hit ? CommitPlugin_logic_free_lineEventStream_fifo_io_pop_payload_mask : 2'b00);
  assign robToPc_valid = FrontendPlugin_allocated_isFireing;
  assign robToPc_robId = FrontendPlugin_allocated_ROB_ID;
  assign robToPc_pc_0 = FrontendPlugin_allocated_PC_0;
  assign robToPc_pc_1 = FrontendPlugin_allocated_PC_1;
  assign commit_robId = CommitPlugin_logic_commit_event_robId;
  assign commit_mask = CommitPlugin_logic_commit_event_mask;
  assign reschedule_valid = CommitPlugin_logic_commit_reschedulePort_valid;
  assign reschedule_payload_robId = CommitPlugin_logic_commit_reschedulePort_payload_robId;
  assign reschedule_payload_robIdNext = CommitPlugin_logic_commit_reschedulePort_payload_robIdNext;
  assign reschedule_payload_trap = CommitPlugin_logic_commit_reschedulePort_payload_trap;
  assign reschedule_payload_cause = CommitPlugin_logic_commit_reschedulePort_payload_cause;
  assign reschedule_payload_tval = CommitPlugin_logic_commit_reschedulePort_payload_tval;
  assign reschedule_payload_reason = CommitPlugin_logic_commit_reschedulePort_payload_reason;
  assign reschedule_payload_skipCommit = CommitPlugin_logic_commit_reschedulePort_payload_skipCommit;
  assign rescheduleReason = CommitPlugin_logic_reschedule_reason;
  assign commit_pc_0 = _zz_commit_pc_0_1[31 : 0];
  assign commit_pc_1 = _zz_commit_pc_0_1[63 : 32];
  assign _zz_CommitDebugFilterPlugin_logic_commits = CommitPlugin_logic_commit_event_mask[0];
  assign _zz_CommitDebugFilterPlugin_logic_commits_1 = CommitPlugin_logic_commit_event_mask[1];
  assign CommitDebugFilterPlugin_logic_commits = ({16'd0,_zz_CommitDebugFilterPlugin_logic_commits_2} <<< 5'd16);
  assign PrivilegedPlugin_logic_defaultTrap_csrPrivilege = EU0_CsrAccessPlugin_setup_onDecodeAddress[9 : 8];
  assign PrivilegedPlugin_logic_defaultTrap_csrReadOnly = (&EU0_CsrAccessPlugin_setup_onDecodeAddress[11 : 10]);
  assign when_PrivilegedPlugin_l165 = ((PrivilegedPlugin_logic_defaultTrap_csrReadOnly && EU0_CsrAccessPlugin_setup_onDecodeWrite) || (PrivilegedPlugin_setup_privilege < PrivilegedPlugin_logic_defaultTrap_csrPrivilege));
  always @(*) begin
    PrivilegedPlugin_logic_machine_mstatus_sd = 1'b0;
    if(when_PrivilegedPlugin_l393) begin
      PrivilegedPlugin_logic_machine_mstatus_sd = 1'b1;
    end
  end

  assign when_PrivilegedPlugin_l393 = (PrivilegedPlugin_logic_machine_mstatus_fs == 2'b11);
  assign PrivilegedPlugin_logic_supervisor_sip_seipOr = (PrivilegedPlugin_logic_supervisor_sip_seipSoft || PrivilegedPlugin_logic_supervisor_sip_seipInput);
  assign PrivilegedPlugin_logic_supervisor_sip_seipMasked = (PrivilegedPlugin_logic_supervisor_sip_seipOr && PrivilegedPlugin_logic_machine_mideleg_se);
  assign PrivilegedPlugin_logic_supervisor_sip_stipMasked = (PrivilegedPlugin_logic_supervisor_sip_stip && PrivilegedPlugin_logic_machine_mideleg_st);
  assign PrivilegedPlugin_logic_supervisor_sip_ssipMasked = (PrivilegedPlugin_logic_supervisor_sip_ssip && PrivilegedPlugin_logic_machine_mideleg_ss);
  assign _zz_when_PrivilegedPlugin_l637 = (PrivilegedPlugin_logic_supervisor_sip_ssip && PrivilegedPlugin_logic_supervisor_sie_ssie);
  assign _zz_when_PrivilegedPlugin_l637_1 = (PrivilegedPlugin_logic_supervisor_sip_stip && PrivilegedPlugin_logic_supervisor_sie_stie);
  assign _zz_when_PrivilegedPlugin_l637_2 = (PrivilegedPlugin_logic_supervisor_sip_seipOr && PrivilegedPlugin_logic_supervisor_sie_seie);
  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_ready = PrivilegedPlugin_logic_reschedule_ready;
    if(when_Stream_l369) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_ready = 1'b1;
    end
  end

  assign when_Stream_l369 = (! PrivilegedPlugin_logic_reschedule_valid);
  assign PrivilegedPlugin_logic_reschedule_valid = PrivilegedPlugin_logic_rescheduleUnbuffered_rValid;
  assign PrivilegedPlugin_logic_reschedule_payload_cause = PrivilegedPlugin_logic_rescheduleUnbuffered_rData_cause;
  assign PrivilegedPlugin_logic_reschedule_payload_epc = PrivilegedPlugin_logic_rescheduleUnbuffered_rData_epc;
  assign PrivilegedPlugin_logic_reschedule_payload_tval = PrivilegedPlugin_logic_rescheduleUnbuffered_rData_tval;
  assign PrivilegedPlugin_logic_reschedule_payload_fromCommit = PrivilegedPlugin_logic_rescheduleUnbuffered_rData_fromCommit;
  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_valid = (CommitPlugin_logic_commit_reschedulePort_valid && CommitPlugin_logic_commit_reschedulePort_payload_trap);
    if(when_PrivilegedPlugin_l585) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_valid = 1'b1;
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_payload_cause = CommitPlugin_logic_commit_reschedulePort_payload_cause;
    if(when_PrivilegedPlugin_l585) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_payload_cause = DecoderPlugin_setup_exceptionPort_payload_cause;
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc = _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_2[31 : 0];
    if(when_PrivilegedPlugin_l585) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc = DecoderPlugin_setup_exceptionPort_payload_epc;
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_rescheduleUnbuffered_payload_tval = CommitPlugin_logic_commit_reschedulePort_payload_tval;
    if(when_PrivilegedPlugin_l585) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_payload_tval = DecoderPlugin_setup_exceptionPort_payload_tval;
    end
  end

  assign PrivilegedPlugin_logic_rescheduleUnbuffered_payload_fromCommit = (CommitPlugin_logic_commit_reschedulePort_valid && CommitPlugin_logic_commit_reschedulePort_payload_trap);
  assign when_PrivilegedPlugin_l585 = (DecoderPlugin_setup_exceptionPort_valid && (! PrivilegedPlugin_logic_rescheduleUnbuffered_payload_fromCommit));
  assign PrivilegedPlugin_logic_targetMachine = 1'b1;
  always @(*) begin
    PrivilegedPlugin_logic_reschedule_ready = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
        PrivilegedPlugin_logic_reschedule_ready = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_branchMissEvent = _zz_PerformanceCounterPlugin_logic_branchMissEvent;
  always @(*) begin
    PerformanceCounterPlugin_logic_commitCount = _zz_PerformanceCounterPlugin_logic_commitCount;
    if(PerformanceCounterPlugin_logic_ignoreNextCommit) begin
      PerformanceCounterPlugin_logic_commitCount = 2'b00;
    end
  end

  assign when_PerformanceCounterPlugin_l65 = (|CommitPlugin_logic_commit_event_mask);
  assign PerformanceCounterPlugin_logic_events_sums_0 = _zz_PerformanceCounterPlugin_logic_events_sums_0;
  assign PerformanceCounterPlugin_logic_events_sums_1 = _zz_PerformanceCounterPlugin_logic_events_sums_1;
  assign PerformanceCounterPlugin_logic_events_sums_2 = _zz_PerformanceCounterPlugin_logic_events_sums_2;
  assign PerformanceCounterPlugin_logic_events_sums_3 = _zz_PerformanceCounterPlugin_logic_events_sums_3;
  always @(*) begin
    _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_1 = 6'h00;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
        if(when_PerformanceCounterPlugin_l201) begin
          case(PerformanceCounterPlugin_logic_fsm_cmd_address)
            3'b001 : begin
              _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_1[5] = 1'b0;
            end
            default : begin
            end
          endcase
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_wantStart = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
        PerformanceCounterPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_fsm_wantKill = 1'b0;
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
        if(!PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
          if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
            PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready = 1'b1;
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_flusherCmd_ready = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
        if(PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
          PerformanceCounterPlugin_logic_fsm_flusherCmd_ready = 1'b1;
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
        PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign ALU0_IntFormatPlugin_logic_stages_0_hits = {ALU0_BranchPlugin_setup_intFormatPort_valid,{ALU0_ShiftPlugin_setup_intFormatPort_valid,ALU0_IntAluPlugin_setup_intFormatPort_valid}};
  assign ALU0_IntFormatPlugin_logic_stages_0_wb_valid = (ALU0_ExecutionUnitBase_pipeline_execute_0_valid && (|ALU0_IntFormatPlugin_logic_stages_0_hits));
  assign ALU0_IntFormatPlugin_logic_stages_0_raw = (((ALU0_IntFormatPlugin_logic_stages_0_hits[0] ? ALU0_IntAluPlugin_setup_intFormatPort_payload : 32'h00000000) | (ALU0_IntFormatPlugin_logic_stages_0_hits[1] ? ALU0_ShiftPlugin_setup_intFormatPort_payload : 32'h00000000)) | (ALU0_IntFormatPlugin_logic_stages_0_hits[2] ? ALU0_BranchPlugin_setup_intFormatPort_payload : 32'h00000000));
  assign ALU0_IntFormatPlugin_logic_stages_0_wb_payload = ALU0_IntFormatPlugin_logic_stages_0_raw;
  always @(*) begin
    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC1_CTRL)
      1'b0 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
      end
      default : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = {ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 12],12'h000};
      end
    endcase
  end

  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  always @(*) begin
    _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL)
      2'b00 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
      end
      2'b01 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = {{20{_zz__zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2[11]}}, _zz__zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2};
      end
      2'b10 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = ALU0_ExecutionUnitBase_pipeline_fetch_0_PC;
      end
      default : begin
      end
    endcase
  end

  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  always @(*) begin
    ALU0_SrcPlugin_logic_addsub_rs2Patched = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
    if(ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT) begin
      ALU0_SrcPlugin_logic_addsub_rs2Patched = (~ ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
    end
    if(ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO) begin
      ALU0_SrcPlugin_logic_addsub_rs2Patched = 32'h00000000;
    end
  end

  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(_zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB) + $signed(_zz_ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1));
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS = ((ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31] == ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31]) ? ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB[31] : (ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED ? ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31] : ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]));
  assign ALU0_IntAluPlugin_setup_intFormatPort_valid = ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_SEL;
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        ALU0_IntAluPlugin_logic_process_bitwise = (ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 & ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        ALU0_IntAluPlugin_logic_process_bitwise = (ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 | ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
      end
      default : begin
        ALU0_IntAluPlugin_logic_process_bitwise = (ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 ^ ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
      end
    endcase
  end

  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_BITWISE : begin
        ALU0_IntAluPlugin_logic_process_result = ALU0_IntAluPlugin_logic_process_bitwise;
      end
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : begin
        ALU0_IntAluPlugin_logic_process_result = _zz_ALU0_IntAluPlugin_logic_process_result;
      end
      default : begin
        ALU0_IntAluPlugin_logic_process_result = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
      end
    endcase
  end

  assign ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_RESULT = ALU0_IntAluPlugin_logic_process_result;
  assign ALU0_IntAluPlugin_setup_intFormatPort_payload = ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_RESULT;
  assign ALU0_ShiftPlugin_setup_intFormatPort_valid = ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SEL;
  assign ALU0_ShiftPlugin_logic_process_amplitude = _zz_ALU0_ShiftPlugin_logic_process_amplitude;
  assign ALU0_ShiftPlugin_logic_process_reversed = (ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT ? _zz_ALU0_ShiftPlugin_logic_process_reversed : ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1);
  assign ALU0_ShiftPlugin_logic_process_shifted = _zz_ALU0_ShiftPlugin_logic_process_shifted[31:0];
  assign ALU0_ShiftPlugin_logic_process_patched = (ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT ? _zz_ALU0_ShiftPlugin_logic_process_patched : ALU0_ShiftPlugin_logic_process_shifted);
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SHIFT_RESULT = ALU0_ShiftPlugin_logic_process_patched;
  assign ALU0_ShiftPlugin_setup_intFormatPort_payload = ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SHIFT_RESULT;
  assign ALU0_BranchPlugin_setup_intFormatPort_valid = ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ = ($signed(ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1) == $signed(ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2));
  assign switch_Misc_l232 = ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[14 : 12];
  always @(*) begin
    casez(switch_Misc_l232)
      3'b000 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ;
      end
      3'b001 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = (! ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ);
      end
      3'b1?1 : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = (! ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS);
      end
      default : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
      end
    endcase
  end

  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1 = 1'b1;
      end
      default : begin
        _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1 = _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
      end
    endcase
  end

  assign ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1;
  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        ALU0_BranchPlugin_logic_process_target_a = ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1;
      end
      default : begin
        ALU0_BranchPlugin_logic_process_target_a = ALU0_ExecutionUnitBase_pipeline_execute_0_PC;
      end
    endcase
  end

  always @(*) begin
    case(ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_JAL : begin
        ALU0_BranchPlugin_logic_process_target_b = {{11{_zz_ALU0_BranchPlugin_logic_process_target_b[20]}}, _zz_ALU0_BranchPlugin_logic_process_target_b};
      end
      BranchPlugin_BranchCtrlEnum_JALR : begin
        ALU0_BranchPlugin_logic_process_target_b = {{20{_zz_ALU0_BranchPlugin_logic_process_target_b_1[11]}}, _zz_ALU0_BranchPlugin_logic_process_target_b_1};
      end
      default : begin
        ALU0_BranchPlugin_logic_process_target_b = {{19{_zz_ALU0_BranchPlugin_logic_process_target_b_2[12]}}, _zz_ALU0_BranchPlugin_logic_process_target_b_2};
      end
    endcase
  end

  always @(*) begin
    ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE = _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE;
    ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE[0] = 1'b0;
  end

  assign ALU0_BranchPlugin_logic_process_slices = (_zz_ALU0_BranchPlugin_logic_process_slices + {1'b0,1'b1});
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE = (ALU0_ExecutionUnitBase_pipeline_execute_0_PC + _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE);
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TARGET = (ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND ? ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE : ALU0_ExecutionUnitBase_pipeline_execute_0_PC_FALSE);
  assign EU0_IntFormatPlugin_logic_stages_0_hits = {EU0_CsrAccessPlugin_setup_intFormatPort_valid,{EU0_DivPlugin_setup_intFormatPort_valid,EU0_MulPlugin_setup_intFormatPort_valid}};
  assign EU0_IntFormatPlugin_logic_stages_0_wb_valid = (EU0_ExecutionUnitBase_pipeline_execute_2_valid && (|EU0_IntFormatPlugin_logic_stages_0_hits));
  assign EU0_IntFormatPlugin_logic_stages_0_raw = (((EU0_IntFormatPlugin_logic_stages_0_hits[0] ? EU0_MulPlugin_setup_intFormatPort_payload : 32'h00000000) | (EU0_IntFormatPlugin_logic_stages_0_hits[1] ? EU0_DivPlugin_setup_intFormatPort_payload : 32'h00000000)) | (EU0_IntFormatPlugin_logic_stages_0_hits[2] ? EU0_CsrAccessPlugin_setup_intFormatPort_payload : 32'h00000000));
  assign EU0_IntFormatPlugin_logic_stages_0_wb_payload = EU0_IntFormatPlugin_logic_stages_0_raw;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
  end

  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(EU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL)
      1'b0 : begin
        _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = {{20{_zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2[11]}}, _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2};
      end
      default : begin
        _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = {{20{_zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2_1[11]}}, _zz__zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2_1};
      end
    endcase
  end

  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  always @(*) begin
    EU0_SrcPlugin_logic_addsub_rs2Patched = EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
    if(EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT) begin
      EU0_SrcPlugin_logic_addsub_rs2Patched = (~ EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO) begin
      EU0_SrcPlugin_logic_addsub_rs2Patched = 32'h00000000;
    end
  end

  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB) + $signed(_zz_EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1));
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS = ((EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31] == EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31]) ? EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB[31] : (EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED ? EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31] : EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]));
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED = EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED = EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT = (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_SIGNED && EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED[31]);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT = (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED && EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED[31]);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED = ((EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT ? (~ EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED) : EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_FORMATED) + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_UNSIGNED);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED = ((EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT ? (~ EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED) : EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED) + _zz_EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_UNSIGNED);
  assign EU0_MulPlugin_setup_intFormatPort_valid = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL;
  assign EU0_MulPlugin_logic_wake_wakeRobsSel = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL;
  assign EU0_MulPlugin_logic_wake_wakeRegFileSel = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1 = {(EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_SIGNED && EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1[31]),EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1};
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2 = {(EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED && EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2[31]),EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2};
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_0 = (EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC1[16 : 0] * EU0_ExecutionUnitBase_pipeline_execute_0_MUL_SRC2[16 : 0]);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3 = _zz_EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0 = 61'h0000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0[33 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_0[33 : 0];
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0[60 : 34] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_3[26 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_1 = 61'h0000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_1[60 : 17] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_1[43 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_2 = 61'h0000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_2[60 : 17] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_2[43 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1 = 3'b000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1[2 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_3[29 : 27];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_1 = 3'b000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_1[2 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_1[46 : 44];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_2 = 3'b000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_2[2 : 0] = EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_2[46 : 44];
  end

  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_3 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0_6);
  assign EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_3 + _zz_EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1_6);
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0 = 66'h00000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0[62 : 0] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_0_adders_0[62 : 0];
  end

  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0_1 = 66'h00000000000000000;
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0_1[65 : 61] = EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_0_adders_1[4 : 0];
  end

  assign EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0 = (_zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0 + _zz_EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0_1);
  assign EU0_MulPlugin_setup_intFormatPort_payload = (EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_HIGH ? EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0[63 : 32] : EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_1_adders_0[31 : 0]);
  assign EU0_DivPlugin_setup_intFormatPort_valid = EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL;
  assign EU0_DivPlugin_logic_wake_wakeRobsSel = EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL;
  assign EU0_DivPlugin_logic_wake_wakeRegFileSel = EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_DIV_REVERT_RESULT = ((EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_REVERT ^ (EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_REVERT && (! EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM))) && (! (((EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_FORMATED == 32'h00000000) && EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED) && (! EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM))));
  assign toplevel_EU0_DivPlugin_logic_div_io_cmd_fire = (EU0_DivPlugin_logic_div_io_cmd_valid && EU0_DivPlugin_logic_div_io_cmd_ready);
  assign when_DivPlugin_l76 = (EU0_ExecutionUnitBase_pipeline_execute_0_ready || EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed);
  assign EU0_DivPlugin_logic_div_io_cmd_valid = ((EU0_ExecutionUnitBase_pipeline_execute_0_valid && EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL) && (! EU0_DivPlugin_logic_feed_cmdSent));
  assign EU0_ExecutionUnitBase_pipeline_execute_0_haltRequest_DivPlugin_l83 = ((EU0_ExecutionUnitBase_pipeline_execute_0_valid && EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL) && (! EU0_DivPlugin_logic_feed_cmdSent));
  assign EU0_ExecutionUnitBase_pipeline_execute_1_haltRequest_DivPlugin_l91 = ((EU0_ExecutionUnitBase_pipeline_execute_1_valid && EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_SEL) && (! EU0_DivPlugin_logic_div_io_rsp_valid));
  assign EU0_DivPlugin_logic_rsp_selected = (EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_REM ? _zz_EU0_DivPlugin_logic_rsp_selected : EU0_DivPlugin_logic_div_io_rsp_payload_result);
  assign _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT = EU0_DivPlugin_logic_rsp_selected;
  assign EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT = _zz_EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT_1[31:0];
  assign EU0_DivPlugin_setup_intFormatPort_payload = EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_DIV_RESULT;
  assign AguPlugin_logic_func3 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[14 : 12];
  assign when_AguPlugin_l89 = (EU0_ExecutionUnitBase_pipeline_execute_0_ready || EU0_ExecutionUnitBase_pipeline_execute_0_isRemoved);
  assign AguPlugin_setup_port_valid = ((EU0_ExecutionUnitBase_pipeline_execute_0_valid && EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SEL) && (! AguPlugin_logic_fired));
  assign AguPlugin_setup_port_payload_address = EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
  assign AguPlugin_setup_port_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  assign AguPlugin_setup_port_payload_robIdMsb = EU0_ExecutionUnitBase_pipeline_execute_0_ROB_MSB;
  assign AguPlugin_setup_port_payload_size = AguPlugin_logic_func3[1 : 0];
  assign AguPlugin_setup_port_payload_sc = EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SC;
  assign AguPlugin_setup_port_payload_amo = EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_AMO;
  assign AguPlugin_setup_port_payload_swap = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[27];
  assign AguPlugin_setup_port_payload_op = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 29];
  assign AguPlugin_setup_port_payload_physicalRd = EU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  assign AguPlugin_setup_port_payload_writeRd = EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD;
  assign AguPlugin_setup_port_payload_aguId = EU0_ExecutionUnitBase_pipeline_execute_0_LSU_ID;
  assign AguPlugin_setup_port_payload_unsigned = AguPlugin_logic_func3[2];
  assign AguPlugin_setup_port_payload_pc = EU0_ExecutionUnitBase_pipeline_execute_0_PC;
  assign AguPlugin_setup_port_payload_lr = EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LR;
  assign AguPlugin_setup_port_payload_load = EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LOAD;
  assign AguPlugin_setup_port_payload_data = EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2;
  assign EnvCallPlugin_setup_reschedule_valid = (EU0_ExecutionUnitBase_pipeline_execute_2_valid && (((((EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA));
  assign EnvCallPlugin_setup_reschedule_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  always @(*) begin
    EnvCallPlugin_setup_reschedule_payload_tval = (EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK ? EU0_ExecutionUnitBase_pipeline_execute_2_PC : 32'h00000000);
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET) begin
      EnvCallPlugin_setup_reschedule_payload_tval[1 : 0] = EnvCallPlugin_logic_xretPriv;
    end
  end

  always @(*) begin
    EnvCallPlugin_setup_reschedule_payload_skipCommit = (EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL);
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET) begin
      if(when_EnvCallPlugin_l95) begin
        EnvCallPlugin_setup_reschedule_payload_skipCommit = 1'b1;
      end
    end
  end

  always @(*) begin
    EnvCallPlugin_setup_reschedule_payload_reason = 8'h02;
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET) begin
      if(when_EnvCallPlugin_l95) begin
        EnvCallPlugin_setup_reschedule_payload_reason = 8'h01;
      end
    end
  end

  always @(*) begin
    EnvCallPlugin_setup_reschedule_payload_cause = 4'bxxxx;
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET) begin
      EnvCallPlugin_setup_reschedule_payload_cause = 4'b1000;
      if(when_EnvCallPlugin_l95) begin
        EnvCallPlugin_setup_reschedule_payload_cause = 4'b0010;
      end
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK) begin
      EnvCallPlugin_setup_reschedule_payload_cause = 4'b0011;
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL) begin
      EnvCallPlugin_setup_reschedule_payload_cause = 4'b1011;
    end
    if(when_EnvCallPlugin_l108) begin
      EnvCallPlugin_setup_reschedule_payload_cause = 4'b1001;
    end
  end

  assign EnvCallPlugin_logic_xretPriv = EU0_ExecutionUnitBase_pipeline_execute_2_Frontend_MICRO_OP[29 : 28];
  assign when_EnvCallPlugin_l95 = (EnvCallPlugin_logic_xretPriv < PrivilegedPlugin_setup_privilege);
  assign when_EnvCallPlugin_l108 = ((EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA) || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA);
  assign EnvCallPlugin_logic_flushes_wantExit = 1'b0;
  always @(*) begin
    EnvCallPlugin_logic_flushes_wantStart = 1'b0;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
        EnvCallPlugin_logic_flushes_wantStart = 1'b1;
      end
    endcase
  end

  assign EnvCallPlugin_logic_flushes_wantKill = 1'b0;
  assign FetchPlugin_stages_0_haltRequest_EnvCallPlugin_l125 = (! (EnvCallPlugin_logic_flushes_stateReg == EnvCallPlugin_logic_flushes_enumDef_IDLE));
  always @(*) begin
    EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_stateReg;
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
        if(EU0_ExecutionUnitBase_pipeline_execute_2_valid) begin
          if(EU0_ExecutionUnitBase_pipeline_execute_2_ready) begin
            if(when_EnvCallPlugin_l135) begin
              EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE;
            end
            if(EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA) begin
              EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH;
            end
          end
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
        if(CommitPlugin_logic_commit_reschedulePort_valid) begin
          EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
        EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT;
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
        if(FetchCachePlugin_setup_invalidatePort_rsp_valid) begin
          EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH;
        end
        if(MmuPlugin_setup_invalidatePort_rsp_valid) begin
          EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_IDLE;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
        EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU;
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
        if(Lsu2Plugin_setup_flushPort_rsp_valid) begin
          EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(EnvCallPlugin_logic_flushes_wantStart) begin
      EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_IDLE;
    end
    if(EnvCallPlugin_logic_flushes_wantKill) begin
      EnvCallPlugin_logic_flushes_stateNext = EnvCallPlugin_logic_flushes_enumDef_BOOT;
    end
  end

  assign when_EnvCallPlugin_l135 = (EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I || EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA);
  assign EU0_CsrAccessPlugin_setup_intFormatPort_valid = EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL;
  assign EU0_CsrAccessPlugin_logic_wake_wakeRobsSel = EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL;
  assign EU0_CsrAccessPlugin_logic_wake_wakeRegFileSel = EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL;
  assign ALU1_IntFormatPlugin_logic_stages_0_hits = {ALU1_BranchPlugin_setup_intFormatPort_valid,{ALU1_ShiftPlugin_setup_intFormatPort_valid,ALU1_IntAluPlugin_setup_intFormatPort_valid}};
  assign ALU1_IntFormatPlugin_logic_stages_0_wb_valid = (ALU1_ExecutionUnitBase_pipeline_execute_0_valid && (|ALU1_IntFormatPlugin_logic_stages_0_hits));
  assign ALU1_IntFormatPlugin_logic_stages_0_raw = (((ALU1_IntFormatPlugin_logic_stages_0_hits[0] ? ALU1_IntAluPlugin_setup_intFormatPort_payload : 32'h00000000) | (ALU1_IntFormatPlugin_logic_stages_0_hits[1] ? ALU1_ShiftPlugin_setup_intFormatPort_payload : 32'h00000000)) | (ALU1_IntFormatPlugin_logic_stages_0_hits[2] ? ALU1_BranchPlugin_setup_intFormatPort_payload : 32'h00000000));
  assign ALU1_IntFormatPlugin_logic_stages_0_wb_payload = ALU1_IntFormatPlugin_logic_stages_0_raw;
  always @(*) begin
    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC1_CTRL)
      1'b0 : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = ALU1_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
      end
      default : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = {ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP[31 : 12],12'h000};
      end
    endcase
  end

  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
  always @(*) begin
    _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL)
      2'b00 : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = ALU1_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
      end
      2'b01 : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = {{20{_zz__zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2[11]}}, _zz__zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2};
      end
      2'b10 : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = ALU1_ExecutionUnitBase_pipeline_fetch_0_PC;
      end
      default : begin
      end
    endcase
  end

  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
  always @(*) begin
    ALU1_SrcPlugin_logic_addsub_rs2Patched = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2;
    if(ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT) begin
      ALU1_SrcPlugin_logic_addsub_rs2Patched = (~ ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
    end
    if(ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO) begin
      ALU1_SrcPlugin_logic_addsub_rs2Patched = 32'h00000000;
    end
  end

  assign ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB = ($signed(_zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB) + $signed(_zz_ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB_1));
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS = ((ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31] == ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31]) ? ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB[31] : (ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED ? ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2[31] : ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1[31]));
  assign ALU1_IntAluPlugin_setup_intFormatPort_valid = ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_SEL;
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        ALU1_IntAluPlugin_logic_process_bitwise = (ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 & ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        ALU1_IntAluPlugin_logic_process_bitwise = (ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 | ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
      end
      default : begin
        ALU1_IntAluPlugin_logic_process_bitwise = (ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 ^ ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2);
      end
    endcase
  end

  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL)
      IntAluPlugin_AluCtrlEnum_BITWISE : begin
        ALU1_IntAluPlugin_logic_process_result = ALU1_IntAluPlugin_logic_process_bitwise;
      end
      IntAluPlugin_AluCtrlEnum_SLT_SLTU : begin
        ALU1_IntAluPlugin_logic_process_result = _zz_ALU1_IntAluPlugin_logic_process_result;
      end
      default : begin
        ALU1_IntAluPlugin_logic_process_result = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ADD_SUB;
      end
    endcase
  end

  assign ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_RESULT = ALU1_IntAluPlugin_logic_process_result;
  assign ALU1_IntAluPlugin_setup_intFormatPort_payload = ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_RESULT;
  assign ALU1_ShiftPlugin_setup_intFormatPort_valid = ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SEL;
  assign ALU1_ShiftPlugin_logic_process_amplitude = _zz_ALU1_ShiftPlugin_logic_process_amplitude;
  assign ALU1_ShiftPlugin_logic_process_reversed = (ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT ? _zz_ALU1_ShiftPlugin_logic_process_reversed : ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1);
  assign ALU1_ShiftPlugin_logic_process_shifted = _zz_ALU1_ShiftPlugin_logic_process_shifted[31:0];
  assign ALU1_ShiftPlugin_logic_process_patched = (ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT ? _zz_ALU1_ShiftPlugin_logic_process_patched : ALU1_ShiftPlugin_logic_process_shifted);
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SHIFT_RESULT = ALU1_ShiftPlugin_logic_process_patched;
  assign ALU1_ShiftPlugin_setup_intFormatPort_payload = ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SHIFT_RESULT;
  assign ALU1_BranchPlugin_setup_intFormatPort_valid = ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ = ($signed(ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1) == $signed(ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2));
  assign switch_Misc_l232_1 = ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[14 : 12];
  always @(*) begin
    casez(switch_Misc_l232_1)
      3'b000 : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ;
      end
      3'b001 : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = (! ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_EQ);
      end
      3'b1?1 : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = (! ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS);
      end
      default : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_LESS;
      end
    endcase
  end

  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1 = 1'b1;
      end
      default : begin
        _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1 = _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
      end
    endcase
  end

  assign ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND = _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND_1;
  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        ALU1_BranchPlugin_logic_process_target_a = ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1;
      end
      default : begin
        ALU1_BranchPlugin_logic_process_target_a = ALU1_ExecutionUnitBase_pipeline_execute_0_PC;
      end
    endcase
  end

  always @(*) begin
    case(ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL)
      BranchPlugin_BranchCtrlEnum_JAL : begin
        ALU1_BranchPlugin_logic_process_target_b = {{11{_zz_ALU1_BranchPlugin_logic_process_target_b[20]}}, _zz_ALU1_BranchPlugin_logic_process_target_b};
      end
      BranchPlugin_BranchCtrlEnum_JALR : begin
        ALU1_BranchPlugin_logic_process_target_b = {{20{_zz_ALU1_BranchPlugin_logic_process_target_b_1[11]}}, _zz_ALU1_BranchPlugin_logic_process_target_b_1};
      end
      default : begin
        ALU1_BranchPlugin_logic_process_target_b = {{19{_zz_ALU1_BranchPlugin_logic_process_target_b_2[12]}}, _zz_ALU1_BranchPlugin_logic_process_target_b_2};
      end
    endcase
  end

  always @(*) begin
    ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TRUE = _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TRUE;
    ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TRUE[0] = 1'b0;
  end

  assign ALU1_BranchPlugin_logic_process_slices = (_zz_ALU1_BranchPlugin_logic_process_slices + {1'b0,1'b1});
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE = (ALU1_ExecutionUnitBase_pipeline_execute_0_PC + _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE);
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TARGET = (ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND ? ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TRUE : ALU1_ExecutionUnitBase_pipeline_execute_0_PC_FALSE);
  assign FrontendPlugin_allocated_haltRequest_FrontendPlugin_l67 = CommitPlugin_logic_reschedule_valid;
  always @(*) begin
    integer_RfTranslationPlugin_logic_impl_io_rollback = CommitPlugin_logic_commit_reschedulePort_valid;
    if(integer_RfTranslationPlugin_logic_init_busy) begin
      integer_RfTranslationPlugin_logic_impl_io_rollback = 1'b1;
    end
  end

  assign integer_RfTranslationPlugin_logic_impl_io_writes_0_valid = (((FrontendPlugin_allocated_isFireing && FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0) && FrontendPlugin_allocated_WRITE_RD_0) && 1'b1);
  assign integer_RfTranslationPlugin_logic_impl_io_writes_1_valid = (((FrontendPlugin_allocated_isFireing && FrontendPlugin_allocated_Frontend_DISPATCH_MASK_1) && FrontendPlugin_allocated_WRITE_RD_1) && 1'b1);
  always @(*) begin
    integer_RfTranslationPlugin_logic_impl_io_commits_0_valid = ((CommitPlugin_logic_commit_event_mask[0] && integer_RfTranslationPlugin_logic_onCommit_writeRd_0) && 1'b1);
    if(integer_RfTranslationPlugin_logic_init_busy) begin
      integer_RfTranslationPlugin_logic_impl_io_commits_0_valid = 1'b1;
    end
  end

  always @(*) begin
    integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_address = integer_RfTranslationPlugin_logic_onCommit_archRd_0;
    if(integer_RfTranslationPlugin_logic_init_busy) begin
      integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_address = integer_RfTranslationPlugin_logic_init_counter[4:0];
    end
  end

  always @(*) begin
    integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_data = integer_RfTranslationPlugin_logic_onCommit_physRd_0;
    if(integer_RfTranslationPlugin_logic_init_busy) begin
      integer_RfTranslationPlugin_logic_impl_io_commits_0_payload_data = 6'h00;
    end
  end

  assign integer_RfTranslationPlugin_logic_impl_io_commits_1_valid = ((CommitPlugin_logic_commit_event_mask[1] && integer_RfTranslationPlugin_logic_onCommit_writeRd_1) && 1'b1);
  assign integer_RfTranslationPlugin_logic_init_busy = (! integer_RfTranslationPlugin_logic_init_counter[5]);
  assign when_RfTranslationPlugin_l193 = 1'b1;
  assign integer_RfTranslationPlugin_logic_impl_io_reads_0_cmd_valid = (FrontendPlugin_allocated_WRITE_RD_0 && when_RfTranslationPlugin_l193);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RD_FREE_0 = 6'bxxxxxx;
    if(when_RfTranslationPlugin_l193) begin
      FrontendPlugin_allocated_PHYS_RD_FREE_0 = integer_RfTranslationPlugin_logic_impl_io_reads_0_rsp_payload;
    end
  end

  assign integer_RfTranslationPlugin_logic_impl_io_reads_1_cmd_valid = (FrontendPlugin_allocated_READ_RS_0_0 && 1'b1);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RS_0_0 = 6'bxxxxxx;
    if(1'b1) begin
      FrontendPlugin_allocated_PHYS_RS_0_0 = integer_RfTranslationPlugin_logic_impl_io_reads_1_rsp_payload;
    end
  end

  assign integer_RfTranslationPlugin_logic_impl_io_reads_2_cmd_valid = (FrontendPlugin_allocated_READ_RS_1_0 && 1'b1);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RS_1_0 = 6'bxxxxxx;
    if(1'b1) begin
      FrontendPlugin_allocated_PHYS_RS_1_0 = integer_RfTranslationPlugin_logic_impl_io_reads_2_rsp_payload;
    end
  end

  assign when_RfTranslationPlugin_l193_1 = 1'b1;
  assign integer_RfTranslationPlugin_logic_impl_io_reads_3_cmd_valid = (FrontendPlugin_allocated_WRITE_RD_1 && when_RfTranslationPlugin_l193_1);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RD_FREE_1 = 6'bxxxxxx;
    if(when_RfTranslationPlugin_l193_1) begin
      FrontendPlugin_allocated_PHYS_RD_FREE_1 = integer_RfTranslationPlugin_logic_impl_io_reads_3_rsp_payload;
    end
    if(when_RfTranslationPlugin_l214) begin
      FrontendPlugin_allocated_PHYS_RD_FREE_1 = FrontendPlugin_allocated_PHYS_RD_0;
    end
  end

  assign integer_RfTranslationPlugin_logic_impl_io_reads_4_cmd_valid = (FrontendPlugin_allocated_READ_RS_0_1 && 1'b1);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RS_0_1 = 6'bxxxxxx;
    if(1'b1) begin
      FrontendPlugin_allocated_PHYS_RS_0_1 = integer_RfTranslationPlugin_logic_impl_io_reads_4_rsp_payload;
    end
    if(when_RfTranslationPlugin_l218) begin
      FrontendPlugin_allocated_PHYS_RS_0_1 = FrontendPlugin_allocated_PHYS_RD_0;
    end
  end

  assign integer_RfTranslationPlugin_logic_impl_io_reads_5_cmd_valid = (FrontendPlugin_allocated_READ_RS_1_1 && 1'b1);
  always @(*) begin
    FrontendPlugin_allocated_PHYS_RS_1_1 = 6'bxxxxxx;
    if(1'b1) begin
      FrontendPlugin_allocated_PHYS_RS_1_1 = integer_RfTranslationPlugin_logic_impl_io_reads_5_rsp_payload;
    end
    if(when_RfTranslationPlugin_l218_1) begin
      FrontendPlugin_allocated_PHYS_RS_1_1 = FrontendPlugin_allocated_PHYS_RD_0;
    end
  end

  assign _zz_when_RfTranslationPlugin_l214 = ((FrontendPlugin_allocated_WRITE_RD_0 && FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0) && 1'b1);
  assign when_RfTranslationPlugin_l214 = ((_zz_when_RfTranslationPlugin_l214 && (FrontendPlugin_allocated_ARCH_RD_0 == FrontendPlugin_allocated_ARCH_RD_1)) && 1'b1);
  assign when_RfTranslationPlugin_l218 = ((_zz_when_RfTranslationPlugin_l214 && (FrontendPlugin_allocated_ARCH_RD_0 == FrontendPlugin_allocated_ARCH_RS_0_1)) && 1'b1);
  assign when_RfTranslationPlugin_l218_1 = ((_zz_when_RfTranslationPlugin_l214 && (FrontendPlugin_allocated_ARCH_RD_0 == FrontendPlugin_allocated_ARCH_RS_1_1)) && 1'b1);
  always @(*) begin
    integer_RfAllocationPlugin_logic_allocator_io_push_0_valid = (((CommitPlugin_logic_free_port_valid && integer_RfAllocationPlugin_logic_push_mask_0) && integer_RfAllocationPlugin_logic_push_writeRd_0) && 1'b1);
    if(when_RfAllocationPlugin_l81) begin
      integer_RfAllocationPlugin_logic_allocator_io_push_0_valid = 1'b0;
    end
    if(integer_RfAllocationPlugin_logic_init_busy) begin
      integer_RfAllocationPlugin_logic_allocator_io_push_0_valid = 1'b1;
    end
  end

  always @(*) begin
    integer_RfAllocationPlugin_logic_allocator_io_push_0_payload = (CommitPlugin_logic_free_port_payload_commited[0] ? integer_RfAllocationPlugin_logic_push_physicalRdOld_0 : integer_RfAllocationPlugin_logic_push_physicalRdNew_0);
    if(integer_RfAllocationPlugin_logic_init_busy) begin
      integer_RfAllocationPlugin_logic_allocator_io_push_0_payload = integer_RfAllocationPlugin_logic_init_counter[5:0];
    end
  end

  assign when_RfAllocationPlugin_l81 = (integer_RfAllocationPlugin_logic_allocator_io_push_0_payload == 6'h00);
  always @(*) begin
    integer_RfAllocationPlugin_logic_allocator_io_push_1_valid = (((CommitPlugin_logic_free_port_valid && integer_RfAllocationPlugin_logic_push_mask_1) && integer_RfAllocationPlugin_logic_push_writeRd_1) && 1'b1);
    if(when_RfAllocationPlugin_l81_1) begin
      integer_RfAllocationPlugin_logic_allocator_io_push_1_valid = 1'b0;
    end
  end

  assign integer_RfAllocationPlugin_logic_allocator_io_push_1_payload = (CommitPlugin_logic_free_port_payload_commited[1] ? integer_RfAllocationPlugin_logic_push_physicalRdOld_1 : integer_RfAllocationPlugin_logic_push_physicalRdNew_1);
  assign when_RfAllocationPlugin_l81_1 = (integer_RfAllocationPlugin_logic_allocator_io_push_1_payload == 6'h00);
  assign integer_RfAllocationPlugin_logic_init_busy = (! integer_RfAllocationPlugin_logic_init_counter[6]);
  assign BranchContextPlugin_logic_onCommit_isBranchCommit_0 = (CommitPlugin_logic_commit_event_mask[0] && BranchContextPlugin_logic_onCommit_isBranch_0);
  assign BranchContextPlugin_logic_onCommit_isBranchCommit_1 = (CommitPlugin_logic_commit_event_mask[1] && BranchContextPlugin_logic_onCommit_isBranch_1);
  assign BranchContextPlugin_logic_onCommit_commitedNext = (BranchContextPlugin_logic_ptr_commited + _zz_BranchContextPlugin_logic_onCommit_commitedNext);
  assign HistoryPlugin_logic_onCommit_valueNext = HistoryPlugin_logic_onCommit_value;
  assign HistoryPlugin_logic_onCommit_whitebox_0 = HistoryPlugin_logic_onCommit_valueNext;
  assign when_HistoryPlugin_l90 = (CommitPlugin_logic_commit_event_mask[0] && HistoryPlugin_logic_onCommit_isConditionalBranch_0);
  assign HistoryPlugin_logic_onCommit_whitebox_1 = HistoryPlugin_logic_onCommit_valueNext_1;
  assign when_HistoryPlugin_l90_1 = (CommitPlugin_logic_commit_event_mask[1] && HistoryPlugin_logic_onCommit_isConditionalBranch_1);
  always @(*) begin
    HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_value;
    if(BtbPlugin_setup_historyPush_flush) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_update_pushes_0_stateNext_1;
    end
    if(FetchCachePlugin_setup_historyJump_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = FetchCachePlugin_setup_historyJump_payload_history;
    end
    if(DecoderPredictionPlugin_setup_historyPush_flush) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_update_pushes_2_stateNext_2;
    end
    if(CommitPlugin_logic_reschedule_reschedulePort_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_update_rescheduleFlush_newHistory;
    end
  end

  assign FetchPlugin_stages_0_BRANCH_HISTORY = HistoryPlugin_logic_onFetch_valueNext;
  assign HistoryPlugin_logic_update_pushes_0_stateNext = HistoryPlugin_logic_update_pushes_0_state;
  assign when_HistoryPlugin_l115 = BtbPlugin_setup_historyPush_mask[0];
  assign HistoryPlugin_logic_update_pushes_2_stateNext = HistoryPlugin_logic_update_pushes_2_state;
  assign when_HistoryPlugin_l115_1 = DecoderPredictionPlugin_setup_historyPush_mask[0];
  assign when_HistoryPlugin_l115_2 = DecoderPredictionPlugin_setup_historyPush_mask[1];
  assign HistoryPlugin_logic_update_rescheduleFlush_instHistory = _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_2[23 : 0];
  assign HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch = _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_2[0];
  assign HistoryPlugin_logic_update_rescheduleFlush_isTaken = _zz_HistoryPlugin_logic_update_rescheduleFlush_isTaken[0];
  assign HistoryPlugin_logic_update_rescheduleFlush_newHistory = (HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch ? {HistoryPlugin_logic_update_rescheduleFlush_instHistory[22 : 0],HistoryPlugin_logic_update_rescheduleFlush_isTaken} : HistoryPlugin_logic_update_rescheduleFlush_instHistory);
  assign DecoderPredictionPlugin_logic_ras_healPush = _zz_DecoderPredictionPlugin_logic_ras_healPush_2[3 : 0];
  assign DecoderPredictionPlugin_logic_ras_healPop = (DecoderPredictionPlugin_logic_ras_healPush - 4'b0001);
  assign DecoderPredictionPlugin_logic_decodePatch_rasPushUsed = 1'b0;
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
            Lsu2Plugin_logic_lq_regs_0_allocation = 1'b1;
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
            Lsu2Plugin_logic_lq_regs_0_allocation = 1'b1;
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315) begin
      Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
            Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b1;
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_103) begin
          Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_103) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_0_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_delete = 1'b0;
    if(when_Lsu2Plugin_l454) begin
      Lsu2Plugin_logic_lq_regs_0_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_16) begin
      Lsu2Plugin_logic_lq_regs_0_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_0_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_103) begin
            Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_103) begin
              Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_103) begin
            Lsu2Plugin_logic_lq_regs_0_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_103) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315 = ((((|(Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_0_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_0_waitOn_sqId)));
  assign when_Lsu2Plugin_l338 = (Lsu2Plugin_logic_lq_regs_0_redoSet || Lsu2Plugin_logic_lq_regs_0_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
            Lsu2Plugin_logic_lq_regs_1_allocation = 1'b1;
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
            Lsu2Plugin_logic_lq_regs_1_allocation = 1'b1;
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_1) begin
      Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
            Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b1;
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_104) begin
          Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_104) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_1_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_delete = 1'b0;
    if(when_Lsu2Plugin_l454_1) begin
      Lsu2Plugin_logic_lq_regs_1_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_17) begin
      Lsu2Plugin_logic_lq_regs_1_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_1_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_104) begin
            Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_104) begin
              Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_104) begin
            Lsu2Plugin_logic_lq_regs_1_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_104) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_1 = ((((|(Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_1_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_1_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_1 = (Lsu2Plugin_logic_lq_regs_1_redoSet || Lsu2Plugin_logic_lq_regs_1_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
            Lsu2Plugin_logic_lq_regs_2_allocation = 1'b1;
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
            Lsu2Plugin_logic_lq_regs_2_allocation = 1'b1;
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_2) begin
      Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
            Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b1;
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_105) begin
          Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_105) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_2_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_delete = 1'b0;
    if(when_Lsu2Plugin_l454_2) begin
      Lsu2Plugin_logic_lq_regs_2_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_18) begin
      Lsu2Plugin_logic_lq_regs_2_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_2_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_105) begin
            Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_105) begin
              Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_105) begin
            Lsu2Plugin_logic_lq_regs_2_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_105) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_2 = ((((|(Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_2_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_2_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_2 = (Lsu2Plugin_logic_lq_regs_2_redoSet || Lsu2Plugin_logic_lq_regs_2_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
            Lsu2Plugin_logic_lq_regs_3_allocation = 1'b1;
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
            Lsu2Plugin_logic_lq_regs_3_allocation = 1'b1;
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_3) begin
      Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
            Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b1;
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_106) begin
          Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_106) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_3_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_delete = 1'b0;
    if(when_Lsu2Plugin_l454_3) begin
      Lsu2Plugin_logic_lq_regs_3_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_19) begin
      Lsu2Plugin_logic_lq_regs_3_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_3_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_106) begin
            Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_106) begin
              Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_106) begin
            Lsu2Plugin_logic_lq_regs_3_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_106) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_3 = ((((|(Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_3_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_3_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_3 = (Lsu2Plugin_logic_lq_regs_3_redoSet || Lsu2Plugin_logic_lq_regs_3_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
            Lsu2Plugin_logic_lq_regs_4_allocation = 1'b1;
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
            Lsu2Plugin_logic_lq_regs_4_allocation = 1'b1;
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_4) begin
      Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
            Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b1;
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_107) begin
          Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_107) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_4_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_delete = 1'b0;
    if(when_Lsu2Plugin_l454_4) begin
      Lsu2Plugin_logic_lq_regs_4_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_20) begin
      Lsu2Plugin_logic_lq_regs_4_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_4_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_107) begin
            Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_107) begin
              Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_107) begin
            Lsu2Plugin_logic_lq_regs_4_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_107) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_4 = ((((|(Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_4_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_4_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_4 = (Lsu2Plugin_logic_lq_regs_4_redoSet || Lsu2Plugin_logic_lq_regs_4_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
            Lsu2Plugin_logic_lq_regs_5_allocation = 1'b1;
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
            Lsu2Plugin_logic_lq_regs_5_allocation = 1'b1;
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_5) begin
      Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
            Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b1;
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_108) begin
          Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_108) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_5_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_delete = 1'b0;
    if(when_Lsu2Plugin_l454_5) begin
      Lsu2Plugin_logic_lq_regs_5_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_21) begin
      Lsu2Plugin_logic_lq_regs_5_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_5_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_108) begin
            Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_108) begin
              Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_108) begin
            Lsu2Plugin_logic_lq_regs_5_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_108) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_5 = ((((|(Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_5_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_5_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_5 = (Lsu2Plugin_logic_lq_regs_5_redoSet || Lsu2Plugin_logic_lq_regs_5_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
            Lsu2Plugin_logic_lq_regs_6_allocation = 1'b1;
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
            Lsu2Plugin_logic_lq_regs_6_allocation = 1'b1;
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_6) begin
      Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
            Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b1;
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_109) begin
          Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_109) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_6_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_delete = 1'b0;
    if(when_Lsu2Plugin_l454_6) begin
      Lsu2Plugin_logic_lq_regs_6_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_22) begin
      Lsu2Plugin_logic_lq_regs_6_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_6_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_109) begin
            Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_109) begin
              Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_109) begin
            Lsu2Plugin_logic_lq_regs_6_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_109) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_6 = ((((|(Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_6_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_6_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_6 = (Lsu2Plugin_logic_lq_regs_6_redoSet || Lsu2Plugin_logic_lq_regs_6_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
            Lsu2Plugin_logic_lq_regs_7_allocation = 1'b1;
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
            Lsu2Plugin_logic_lq_regs_7_allocation = 1'b1;
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_7) begin
      Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
            Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b1;
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_110) begin
          Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_110) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_7_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_delete = 1'b0;
    if(when_Lsu2Plugin_l454_7) begin
      Lsu2Plugin_logic_lq_regs_7_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_23) begin
      Lsu2Plugin_logic_lq_regs_7_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_7_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_110) begin
            Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_110) begin
              Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_110) begin
            Lsu2Plugin_logic_lq_regs_7_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_110) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_7 = ((((|(Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_7_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_7_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_7 = (Lsu2Plugin_logic_lq_regs_7_redoSet || Lsu2Plugin_logic_lq_regs_7_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_8_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
            Lsu2Plugin_logic_lq_regs_8_allocation = 1'b1;
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
            Lsu2Plugin_logic_lq_regs_8_allocation = 1'b1;
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_8_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_8) begin
      Lsu2Plugin_logic_lq_regs_8_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
            Lsu2Plugin_logic_lq_regs_8_redoSet = 1'b1;
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_111) begin
          Lsu2Plugin_logic_lq_regs_8_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_111) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_8_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_8_delete = 1'b0;
    if(when_Lsu2Plugin_l454_8) begin
      Lsu2Plugin_logic_lq_regs_8_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_24) begin
      Lsu2Plugin_logic_lq_regs_8_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_8_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_111) begin
            Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_111) begin
              Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_8_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_111) begin
            Lsu2Plugin_logic_lq_regs_8_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_111) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_8 = ((((|(Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_8_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_8_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_8_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_8 = (Lsu2Plugin_logic_lq_regs_8_redoSet || Lsu2Plugin_logic_lq_regs_8_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_9_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
            Lsu2Plugin_logic_lq_regs_9_allocation = 1'b1;
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
            Lsu2Plugin_logic_lq_regs_9_allocation = 1'b1;
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_9_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_9) begin
      Lsu2Plugin_logic_lq_regs_9_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
            Lsu2Plugin_logic_lq_regs_9_redoSet = 1'b1;
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_112) begin
          Lsu2Plugin_logic_lq_regs_9_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_112) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_9_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_9_delete = 1'b0;
    if(when_Lsu2Plugin_l454_9) begin
      Lsu2Plugin_logic_lq_regs_9_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_25) begin
      Lsu2Plugin_logic_lq_regs_9_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_9_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_112) begin
            Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_112) begin
              Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_9_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_112) begin
            Lsu2Plugin_logic_lq_regs_9_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_112) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_9 = ((((|(Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_9_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_9_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_9_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_9 = (Lsu2Plugin_logic_lq_regs_9_redoSet || Lsu2Plugin_logic_lq_regs_9_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_10_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
            Lsu2Plugin_logic_lq_regs_10_allocation = 1'b1;
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
            Lsu2Plugin_logic_lq_regs_10_allocation = 1'b1;
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_10_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_10) begin
      Lsu2Plugin_logic_lq_regs_10_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
            Lsu2Plugin_logic_lq_regs_10_redoSet = 1'b1;
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_113) begin
          Lsu2Plugin_logic_lq_regs_10_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_113) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_10_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_10_delete = 1'b0;
    if(when_Lsu2Plugin_l454_10) begin
      Lsu2Plugin_logic_lq_regs_10_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_26) begin
      Lsu2Plugin_logic_lq_regs_10_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_10_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_113) begin
            Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_113) begin
              Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_10_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_113) begin
            Lsu2Plugin_logic_lq_regs_10_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_113) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_10 = ((((|(Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_10_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_10_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_10_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_10 = (Lsu2Plugin_logic_lq_regs_10_redoSet || Lsu2Plugin_logic_lq_regs_10_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_11_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
            Lsu2Plugin_logic_lq_regs_11_allocation = 1'b1;
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
            Lsu2Plugin_logic_lq_regs_11_allocation = 1'b1;
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_11_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_11) begin
      Lsu2Plugin_logic_lq_regs_11_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
            Lsu2Plugin_logic_lq_regs_11_redoSet = 1'b1;
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_114) begin
          Lsu2Plugin_logic_lq_regs_11_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_114) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_11_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_11_delete = 1'b0;
    if(when_Lsu2Plugin_l454_11) begin
      Lsu2Plugin_logic_lq_regs_11_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_27) begin
      Lsu2Plugin_logic_lq_regs_11_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_11_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_114) begin
            Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_114) begin
              Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_11_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_114) begin
            Lsu2Plugin_logic_lq_regs_11_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_114) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_11 = ((((|(Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_11_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_11_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_11_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_11 = (Lsu2Plugin_logic_lq_regs_11_redoSet || Lsu2Plugin_logic_lq_regs_11_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_12_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
            Lsu2Plugin_logic_lq_regs_12_allocation = 1'b1;
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
            Lsu2Plugin_logic_lq_regs_12_allocation = 1'b1;
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_12_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_12) begin
      Lsu2Plugin_logic_lq_regs_12_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
            Lsu2Plugin_logic_lq_regs_12_redoSet = 1'b1;
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_115) begin
          Lsu2Plugin_logic_lq_regs_12_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_115) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_12_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_12_delete = 1'b0;
    if(when_Lsu2Plugin_l454_12) begin
      Lsu2Plugin_logic_lq_regs_12_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_28) begin
      Lsu2Plugin_logic_lq_regs_12_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_12_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_115) begin
            Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_115) begin
              Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_12_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_115) begin
            Lsu2Plugin_logic_lq_regs_12_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_115) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_12 = ((((|(Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_12_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_12_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_12_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_12 = (Lsu2Plugin_logic_lq_regs_12_redoSet || Lsu2Plugin_logic_lq_regs_12_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_13_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
            Lsu2Plugin_logic_lq_regs_13_allocation = 1'b1;
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
            Lsu2Plugin_logic_lq_regs_13_allocation = 1'b1;
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_13_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_13) begin
      Lsu2Plugin_logic_lq_regs_13_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
            Lsu2Plugin_logic_lq_regs_13_redoSet = 1'b1;
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_116) begin
          Lsu2Plugin_logic_lq_regs_13_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_116) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_13_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_13_delete = 1'b0;
    if(when_Lsu2Plugin_l454_13) begin
      Lsu2Plugin_logic_lq_regs_13_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_29) begin
      Lsu2Plugin_logic_lq_regs_13_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_13_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_116) begin
            Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_116) begin
              Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_13_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_116) begin
            Lsu2Plugin_logic_lq_regs_13_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_116) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_13 = ((((|(Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_13_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_13_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_13_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_13 = (Lsu2Plugin_logic_lq_regs_13_redoSet || Lsu2Plugin_logic_lq_regs_13_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_14_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
            Lsu2Plugin_logic_lq_regs_14_allocation = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
            Lsu2Plugin_logic_lq_regs_14_allocation = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_14_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_14) begin
      Lsu2Plugin_logic_lq_regs_14_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
            Lsu2Plugin_logic_lq_regs_14_redoSet = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_117) begin
          Lsu2Plugin_logic_lq_regs_14_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_117) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_14_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_14_delete = 1'b0;
    if(when_Lsu2Plugin_l454_14) begin
      Lsu2Plugin_logic_lq_regs_14_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_30) begin
      Lsu2Plugin_logic_lq_regs_14_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_14_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_117) begin
            Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_117) begin
              Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_14_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_117) begin
            Lsu2Plugin_logic_lq_regs_14_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_117) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_14 = ((((|(Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_14_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_14_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_14_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_14 = (Lsu2Plugin_logic_lq_regs_14_redoSet || Lsu2Plugin_logic_lq_regs_14_delete);
  always @(*) begin
    Lsu2Plugin_logic_lq_regs_15_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
            Lsu2Plugin_logic_lq_regs_15_allocation = 1'b1;
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_LQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
            Lsu2Plugin_logic_lq_regs_15_allocation = 1'b1;
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_15_redoSet = 1'b0;
    if(when_Lsu2Plugin_l315_15) begin
      Lsu2Plugin_logic_lq_regs_15_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_2)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
            Lsu2Plugin_logic_lq_regs_15_redoSet = 1'b1;
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_118) begin
          Lsu2Plugin_logic_lq_regs_15_redoSet = 1'b1;
        end
      end
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_118) begin
            if(when_Lsu2Plugin_l1314) begin
              Lsu2Plugin_logic_lq_regs_15_redoSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_15_delete = 1'b0;
    if(when_Lsu2Plugin_l454_15) begin
      Lsu2Plugin_logic_lq_regs_15_delete = 1'b1;
    end
    if(when_Lsu2Plugin_l454_31) begin
      Lsu2Plugin_logic_lq_regs_15_delete = 1'b1;
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_regs_15_delete = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefillSet = 2'b00;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          if(_zz_118) begin
            Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefillSet = Lsu2Plugin_logic_sharedPip_ctrl_refillMask;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_118) begin
              Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_15_waitOn_sqWritebackSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_118) begin
            Lsu2Plugin_logic_lq_regs_15_waitOn_sqWritebackSet = 1'b1;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeedSet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_118) begin
            if(when_Lsu2Plugin_l1313) begin
              Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeedSet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l315_15 = ((((|(Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefill & DataCachePlugin_setup_refillCompletions)) || (Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake)) || ((Lsu2Plugin_logic_lq_regs_15_waitOn_sqWriteback && Lsu2Plugin_logic_sqWritebackEvent_valid) && (Lsu2Plugin_logic_sqWritebackEvent_payload == Lsu2Plugin_logic_lq_regs_15_waitOn_sqId))) || ((Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeed && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_lq_regs_15_waitOn_sqId)));
  assign when_Lsu2Plugin_l338_15 = (Lsu2Plugin_logic_lq_regs_15_redoSet || Lsu2Plugin_logic_lq_regs_15_delete);
  assign Lsu2Plugin_logic_lq_ptr_allocReal = Lsu2Plugin_logic_lq_ptr_alloc[3 : 0];
  assign Lsu2Plugin_logic_lq_ptr_freeReal = Lsu2Plugin_logic_lq_ptr_free[3 : 0];
  assign when_UInt_l120 = (|Lsu2Plugin_logic_lq_tracker_freeNext[4 : 2]);
  always @(*) begin
    if(when_UInt_l120) begin
      _zz_Lsu2Plugin_logic_lq_tracker_freeReduced = 2'b11;
    end else begin
      _zz_Lsu2Plugin_logic_lq_tracker_freeReduced = Lsu2Plugin_logic_lq_tracker_freeNext[1 : 0];
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_tracker_freeNext = (_zz_Lsu2Plugin_logic_lq_tracker_freeNext - _zz_Lsu2Plugin_logic_lq_tracker_freeNext_2);
    if(Lsu2Plugin_logic_lq_tracker_clear) begin
      Lsu2Plugin_logic_lq_tracker_freeNext = 5'h10;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_tracker_clear = 1'b0;
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lq_tracker_clear = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_lq_onCommit_lqCommits_0 = (CommitPlugin_logic_commit_event_mask[0] && Lsu2Plugin_logic_lq_onCommit_lqAlloc_0);
  assign Lsu2Plugin_logic_lq_onCommit_lqCommits_1 = (CommitPlugin_logic_commit_event_mask[1] && Lsu2Plugin_logic_lq_onCommit_lqAlloc_1);
  assign Lsu2Plugin_logic_lq_onCommit_lqCommitCount = _zz_Lsu2Plugin_logic_lq_onCommit_lqCommitCount;
  assign Lsu2Plugin_logic_lq_onCommit_free = Lsu2Plugin_logic_lq_ptr_free;
  assign Lsu2Plugin_logic_lq_onCommit_priority = Lsu2Plugin_logic_lq_ptr_priority;
  assign when_Lsu2Plugin_l454 = ((_zz_when_Lsu2Plugin_l454 == 4'b0000) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_1 = ((_zz_when_Lsu2Plugin_l454_1 == 4'b0001) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_2 = ((_zz_when_Lsu2Plugin_l454_2 == 4'b0010) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_3 = ((_zz_when_Lsu2Plugin_l454_3 == 4'b0011) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_4 = ((_zz_when_Lsu2Plugin_l454_4 == 4'b0100) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_5 = ((_zz_when_Lsu2Plugin_l454_5 == 4'b0101) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_6 = ((_zz_when_Lsu2Plugin_l454_6 == 4'b0110) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_7 = ((_zz_when_Lsu2Plugin_l454_7 == 4'b0111) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_8 = ((_zz_when_Lsu2Plugin_l454_8 == 4'b1000) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_9 = ((_zz_when_Lsu2Plugin_l454_9 == 4'b1001) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_10 = ((_zz_when_Lsu2Plugin_l454_10 == 4'b1010) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_11 = ((_zz_when_Lsu2Plugin_l454_11 == 4'b1011) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_12 = ((_zz_when_Lsu2Plugin_l454_12 == 4'b1100) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_13 = ((_zz_when_Lsu2Plugin_l454_13 == 4'b1101) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_14 = ((_zz_when_Lsu2Plugin_l454_14 == 4'b1110) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_15 = ((_zz_when_Lsu2Plugin_l454_15 == 4'b1111) && Lsu2Plugin_logic_lq_onCommit_lqCommits_0);
  assign when_Lsu2Plugin_l454_16 = ((_zz_when_Lsu2Plugin_l454_16 == 4'b0000) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_17 = ((_zz_when_Lsu2Plugin_l454_17 == 4'b0001) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_18 = ((_zz_when_Lsu2Plugin_l454_18 == 4'b0010) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_19 = ((_zz_when_Lsu2Plugin_l454_19 == 4'b0011) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_20 = ((_zz_when_Lsu2Plugin_l454_20 == 4'b0100) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_21 = ((_zz_when_Lsu2Plugin_l454_21 == 4'b0101) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_22 = ((_zz_when_Lsu2Plugin_l454_22 == 4'b0110) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_23 = ((_zz_when_Lsu2Plugin_l454_23 == 4'b0111) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_24 = ((_zz_when_Lsu2Plugin_l454_24 == 4'b1000) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_25 = ((_zz_when_Lsu2Plugin_l454_25 == 4'b1001) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_26 = ((_zz_when_Lsu2Plugin_l454_26 == 4'b1010) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_27 = ((_zz_when_Lsu2Plugin_l454_27 == 4'b1011) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_28 = ((_zz_when_Lsu2Plugin_l454_28 == 4'b1100) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_29 = ((_zz_when_Lsu2Plugin_l454_29 == 4'b1101) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_30 = ((_zz_when_Lsu2Plugin_l454_30 == 4'b1110) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign when_Lsu2Plugin_l454_31 = ((_zz_when_Lsu2Plugin_l454_31 == 4'b1111) && Lsu2Plugin_logic_lq_onCommit_lqCommits_1);
  assign Lsu2Plugin_logic_lq_tracker_add = Lsu2Plugin_logic_lq_onCommit_lqCommitCount;
  always @(*) begin
    Lsu2Plugin_logic_lq_reservation_kill = 1'b0;
    if(DataCachePlugin_setup_writebackBusy) begin
      Lsu2Plugin_logic_lq_reservation_kill = 1'b1;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
        if(when_Lsu2Plugin_l1715) begin
          Lsu2Plugin_logic_lq_reservation_kill = 1'b1;
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  assign when_Lsu2Plugin_l484 = Lsu2Plugin_logic_lq_reservation_counter[6];
  assign Lsu2Plugin_logic_lq_hazardPrediction_hazard = 1'b0;
  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_valid = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_VALID;
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_valid = 1'b1;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address = 7'bxxxxxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC[8 : 2];
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC[8 : 2];
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'bxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE + _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score);
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'b111;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag = 16'bxxxxxxxxxxxxxxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC[24 : 9];
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC[24 : 9];
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta = 4'bxxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_DELTA;
          end else begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta = _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta[3:0];
            end
          end
        end
      endcase
    end
  end

  assign _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score = {Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_delta,{Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_tag,Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_score}};
  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_valid = (Lsu2Plugin_logic_lq_hazardPrediction_write_valid && (! Lsu2Plugin_logic_lq_hazardPrediction_hazard));
  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_address = Lsu2Plugin_logic_lq_hazardPrediction_write_payload_address;
  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_score = Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score;
  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_tag = Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_tag;
  assign Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_data_delta = Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_delta;
  assign _zz_when_MultiportRam_l362_2 = Lsu2Plugin_logic_lq_hazardPrediction_write_takeWhen_payload_address;
  assign Lsu2Plugin_logic_lq_hitPrediction_hazard = 1'b0;
  assign _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter = Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_data_counter;
  assign Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_valid = (Lsu2Plugin_logic_lq_hitPrediction_write_valid && (! Lsu2Plugin_logic_lq_hitPrediction_hazard));
  assign Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_address = Lsu2Plugin_logic_lq_hitPrediction_write_payload_address;
  assign Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_data_counter = Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter;
  assign _zz_when_MultiportRam_l362_3 = Lsu2Plugin_logic_lq_hitPrediction_write_takeWhen_payload_address;
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
            Lsu2Plugin_logic_sq_regs_0_allocation = 1'b1;
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
            Lsu2Plugin_logic_sq_regs_0_allocation = 1'b1;
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369) begin
      Lsu2Plugin_logic_sq_regs_0_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
            Lsu2Plugin_logic_sq_regs_0_redoSet = 1'b1;
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_119) begin
          Lsu2Plugin_logic_sq_regs_0_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524) begin
        Lsu2Plugin_logic_sq_regs_0_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909) begin
        Lsu2Plugin_logic_sq_regs_0_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_commitedNext = Lsu2Plugin_logic_sq_regs_0_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[0]) begin
        Lsu2Plugin_logic_sq_regs_0_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[0]) begin
        Lsu2Plugin_logic_sq_regs_0_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_119) begin
              Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369 = (Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385 = (Lsu2Plugin_logic_sq_regs_0_redoSet || Lsu2Plugin_logic_sq_regs_0_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
            Lsu2Plugin_logic_sq_regs_1_allocation = 1'b1;
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
            Lsu2Plugin_logic_sq_regs_1_allocation = 1'b1;
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_1) begin
      Lsu2Plugin_logic_sq_regs_1_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
            Lsu2Plugin_logic_sq_regs_1_redoSet = 1'b1;
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_120) begin
          Lsu2Plugin_logic_sq_regs_1_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_1) begin
        Lsu2Plugin_logic_sq_regs_1_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_1) begin
        Lsu2Plugin_logic_sq_regs_1_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_commitedNext = Lsu2Plugin_logic_sq_regs_1_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[1]) begin
        Lsu2Plugin_logic_sq_regs_1_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[1]) begin
        Lsu2Plugin_logic_sq_regs_1_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_120) begin
              Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_1 = (Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_1 = (Lsu2Plugin_logic_sq_regs_1_redoSet || Lsu2Plugin_logic_sq_regs_1_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
            Lsu2Plugin_logic_sq_regs_2_allocation = 1'b1;
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
            Lsu2Plugin_logic_sq_regs_2_allocation = 1'b1;
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_2) begin
      Lsu2Plugin_logic_sq_regs_2_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
            Lsu2Plugin_logic_sq_regs_2_redoSet = 1'b1;
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_121) begin
          Lsu2Plugin_logic_sq_regs_2_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_2) begin
        Lsu2Plugin_logic_sq_regs_2_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_2) begin
        Lsu2Plugin_logic_sq_regs_2_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_commitedNext = Lsu2Plugin_logic_sq_regs_2_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[2]) begin
        Lsu2Plugin_logic_sq_regs_2_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[2]) begin
        Lsu2Plugin_logic_sq_regs_2_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_121) begin
              Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_2 = (Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_2 = (Lsu2Plugin_logic_sq_regs_2_redoSet || Lsu2Plugin_logic_sq_regs_2_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
            Lsu2Plugin_logic_sq_regs_3_allocation = 1'b1;
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
            Lsu2Plugin_logic_sq_regs_3_allocation = 1'b1;
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_3) begin
      Lsu2Plugin_logic_sq_regs_3_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
            Lsu2Plugin_logic_sq_regs_3_redoSet = 1'b1;
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_122) begin
          Lsu2Plugin_logic_sq_regs_3_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_3) begin
        Lsu2Plugin_logic_sq_regs_3_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_3) begin
        Lsu2Plugin_logic_sq_regs_3_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_commitedNext = Lsu2Plugin_logic_sq_regs_3_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[3]) begin
        Lsu2Plugin_logic_sq_regs_3_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[3]) begin
        Lsu2Plugin_logic_sq_regs_3_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_122) begin
              Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_3 = (Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_3 = (Lsu2Plugin_logic_sq_regs_3_redoSet || Lsu2Plugin_logic_sq_regs_3_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
            Lsu2Plugin_logic_sq_regs_4_allocation = 1'b1;
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
            Lsu2Plugin_logic_sq_regs_4_allocation = 1'b1;
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_4) begin
      Lsu2Plugin_logic_sq_regs_4_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
            Lsu2Plugin_logic_sq_regs_4_redoSet = 1'b1;
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_123) begin
          Lsu2Plugin_logic_sq_regs_4_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_4) begin
        Lsu2Plugin_logic_sq_regs_4_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_4) begin
        Lsu2Plugin_logic_sq_regs_4_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_commitedNext = Lsu2Plugin_logic_sq_regs_4_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[4]) begin
        Lsu2Plugin_logic_sq_regs_4_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[4]) begin
        Lsu2Plugin_logic_sq_regs_4_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_123) begin
              Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_4 = (Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_4 = (Lsu2Plugin_logic_sq_regs_4_redoSet || Lsu2Plugin_logic_sq_regs_4_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
            Lsu2Plugin_logic_sq_regs_5_allocation = 1'b1;
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
            Lsu2Plugin_logic_sq_regs_5_allocation = 1'b1;
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_5) begin
      Lsu2Plugin_logic_sq_regs_5_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
            Lsu2Plugin_logic_sq_regs_5_redoSet = 1'b1;
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_124) begin
          Lsu2Plugin_logic_sq_regs_5_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_5) begin
        Lsu2Plugin_logic_sq_regs_5_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_5) begin
        Lsu2Plugin_logic_sq_regs_5_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_commitedNext = Lsu2Plugin_logic_sq_regs_5_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[5]) begin
        Lsu2Plugin_logic_sq_regs_5_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[5]) begin
        Lsu2Plugin_logic_sq_regs_5_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_124) begin
              Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_5 = (Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_5 = (Lsu2Plugin_logic_sq_regs_5_redoSet || Lsu2Plugin_logic_sq_regs_5_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
            Lsu2Plugin_logic_sq_regs_6_allocation = 1'b1;
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
            Lsu2Plugin_logic_sq_regs_6_allocation = 1'b1;
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_6) begin
      Lsu2Plugin_logic_sq_regs_6_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
            Lsu2Plugin_logic_sq_regs_6_redoSet = 1'b1;
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_125) begin
          Lsu2Plugin_logic_sq_regs_6_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_6) begin
        Lsu2Plugin_logic_sq_regs_6_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_6) begin
        Lsu2Plugin_logic_sq_regs_6_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_commitedNext = Lsu2Plugin_logic_sq_regs_6_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[6]) begin
        Lsu2Plugin_logic_sq_regs_6_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[6]) begin
        Lsu2Plugin_logic_sq_regs_6_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_125) begin
              Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_6 = (Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_6 = (Lsu2Plugin_logic_sq_regs_6_redoSet || Lsu2Plugin_logic_sq_regs_6_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
            Lsu2Plugin_logic_sq_regs_7_allocation = 1'b1;
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
            Lsu2Plugin_logic_sq_regs_7_allocation = 1'b1;
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_7) begin
      Lsu2Plugin_logic_sq_regs_7_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
            Lsu2Plugin_logic_sq_regs_7_redoSet = 1'b1;
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_126) begin
          Lsu2Plugin_logic_sq_regs_7_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_7) begin
        Lsu2Plugin_logic_sq_regs_7_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_7) begin
        Lsu2Plugin_logic_sq_regs_7_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_commitedNext = Lsu2Plugin_logic_sq_regs_7_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[7]) begin
        Lsu2Plugin_logic_sq_regs_7_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[7]) begin
        Lsu2Plugin_logic_sq_regs_7_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_126) begin
              Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_7 = (Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_7 = (Lsu2Plugin_logic_sq_regs_7_redoSet || Lsu2Plugin_logic_sq_regs_7_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_8_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
            Lsu2Plugin_logic_sq_regs_8_allocation = 1'b1;
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
            Lsu2Plugin_logic_sq_regs_8_allocation = 1'b1;
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_8_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_8) begin
      Lsu2Plugin_logic_sq_regs_8_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
            Lsu2Plugin_logic_sq_regs_8_redoSet = 1'b1;
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_127) begin
          Lsu2Plugin_logic_sq_regs_8_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_8_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_8) begin
        Lsu2Plugin_logic_sq_regs_8_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_8) begin
        Lsu2Plugin_logic_sq_regs_8_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_8_commitedNext = Lsu2Plugin_logic_sq_regs_8_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[8]) begin
        Lsu2Plugin_logic_sq_regs_8_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[8]) begin
        Lsu2Plugin_logic_sq_regs_8_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_127) begin
              Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_8 = (Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_8 = (Lsu2Plugin_logic_sq_regs_8_redoSet || Lsu2Plugin_logic_sq_regs_8_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_9_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
            Lsu2Plugin_logic_sq_regs_9_allocation = 1'b1;
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
            Lsu2Plugin_logic_sq_regs_9_allocation = 1'b1;
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_9_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_9) begin
      Lsu2Plugin_logic_sq_regs_9_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
            Lsu2Plugin_logic_sq_regs_9_redoSet = 1'b1;
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_128) begin
          Lsu2Plugin_logic_sq_regs_9_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_9_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_9) begin
        Lsu2Plugin_logic_sq_regs_9_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_9) begin
        Lsu2Plugin_logic_sq_regs_9_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_9_commitedNext = Lsu2Plugin_logic_sq_regs_9_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[9]) begin
        Lsu2Plugin_logic_sq_regs_9_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[9]) begin
        Lsu2Plugin_logic_sq_regs_9_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_128) begin
              Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_9 = (Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_9 = (Lsu2Plugin_logic_sq_regs_9_redoSet || Lsu2Plugin_logic_sq_regs_9_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_10_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
            Lsu2Plugin_logic_sq_regs_10_allocation = 1'b1;
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
            Lsu2Plugin_logic_sq_regs_10_allocation = 1'b1;
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_10_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_10) begin
      Lsu2Plugin_logic_sq_regs_10_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
            Lsu2Plugin_logic_sq_regs_10_redoSet = 1'b1;
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_129) begin
          Lsu2Plugin_logic_sq_regs_10_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_10_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_10) begin
        Lsu2Plugin_logic_sq_regs_10_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_10) begin
        Lsu2Plugin_logic_sq_regs_10_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_10_commitedNext = Lsu2Plugin_logic_sq_regs_10_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[10]) begin
        Lsu2Plugin_logic_sq_regs_10_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[10]) begin
        Lsu2Plugin_logic_sq_regs_10_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_129) begin
              Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_10 = (Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_10 = (Lsu2Plugin_logic_sq_regs_10_redoSet || Lsu2Plugin_logic_sq_regs_10_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_11_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
            Lsu2Plugin_logic_sq_regs_11_allocation = 1'b1;
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
            Lsu2Plugin_logic_sq_regs_11_allocation = 1'b1;
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_11_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_11) begin
      Lsu2Plugin_logic_sq_regs_11_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
            Lsu2Plugin_logic_sq_regs_11_redoSet = 1'b1;
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_130) begin
          Lsu2Plugin_logic_sq_regs_11_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_11_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_11) begin
        Lsu2Plugin_logic_sq_regs_11_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_11) begin
        Lsu2Plugin_logic_sq_regs_11_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_11_commitedNext = Lsu2Plugin_logic_sq_regs_11_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[11]) begin
        Lsu2Plugin_logic_sq_regs_11_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[11]) begin
        Lsu2Plugin_logic_sq_regs_11_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_130) begin
              Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_11 = (Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_11 = (Lsu2Plugin_logic_sq_regs_11_redoSet || Lsu2Plugin_logic_sq_regs_11_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_12_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
            Lsu2Plugin_logic_sq_regs_12_allocation = 1'b1;
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
            Lsu2Plugin_logic_sq_regs_12_allocation = 1'b1;
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_12_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_12) begin
      Lsu2Plugin_logic_sq_regs_12_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
            Lsu2Plugin_logic_sq_regs_12_redoSet = 1'b1;
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_131) begin
          Lsu2Plugin_logic_sq_regs_12_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_12_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_12) begin
        Lsu2Plugin_logic_sq_regs_12_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_12) begin
        Lsu2Plugin_logic_sq_regs_12_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_12_commitedNext = Lsu2Plugin_logic_sq_regs_12_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[12]) begin
        Lsu2Plugin_logic_sq_regs_12_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[12]) begin
        Lsu2Plugin_logic_sq_regs_12_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_131) begin
              Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_12 = (Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_12 = (Lsu2Plugin_logic_sq_regs_12_redoSet || Lsu2Plugin_logic_sq_regs_12_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_13_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
            Lsu2Plugin_logic_sq_regs_13_allocation = 1'b1;
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
            Lsu2Plugin_logic_sq_regs_13_allocation = 1'b1;
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_13_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_13) begin
      Lsu2Plugin_logic_sq_regs_13_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
            Lsu2Plugin_logic_sq_regs_13_redoSet = 1'b1;
          end
          4'b1110 : begin
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_132) begin
          Lsu2Plugin_logic_sq_regs_13_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_13_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_13) begin
        Lsu2Plugin_logic_sq_regs_13_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_13) begin
        Lsu2Plugin_logic_sq_regs_13_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_13_commitedNext = Lsu2Plugin_logic_sq_regs_13_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[13]) begin
        Lsu2Plugin_logic_sq_regs_13_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[13]) begin
        Lsu2Plugin_logic_sq_regs_13_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_132) begin
              Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_13 = (Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_13 = (Lsu2Plugin_logic_sq_regs_13_redoSet || Lsu2Plugin_logic_sq_regs_13_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_14_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
            Lsu2Plugin_logic_sq_regs_14_allocation = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
            Lsu2Plugin_logic_sq_regs_14_allocation = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_14_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_14) begin
      Lsu2Plugin_logic_sq_regs_14_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
            Lsu2Plugin_logic_sq_regs_14_redoSet = 1'b1;
          end
          default : begin
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_133) begin
          Lsu2Plugin_logic_sq_regs_14_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_14_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_14) begin
        Lsu2Plugin_logic_sq_regs_14_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_14) begin
        Lsu2Plugin_logic_sq_regs_14_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_14_commitedNext = Lsu2Plugin_logic_sq_regs_14_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[14]) begin
        Lsu2Plugin_logic_sq_regs_14_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[14]) begin
        Lsu2Plugin_logic_sq_regs_14_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_133) begin
              Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_14 = (Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_14 = (Lsu2Plugin_logic_sq_regs_14_redoSet || Lsu2Plugin_logic_sq_regs_14_delete);
  always @(*) begin
    Lsu2Plugin_logic_sq_regs_15_allocation = 1'b0;
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_0)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
            Lsu2Plugin_logic_sq_regs_15_allocation = 1'b1;
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      if(FrontendPlugin_dispatch_isFireing) begin
        case(FrontendPlugin_dispatch_SQ_ID_1)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
            Lsu2Plugin_logic_sq_regs_15_allocation = 1'b1;
          end
        endcase
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_15_redoSet = 1'b0;
    if(when_Lsu2Plugin_l369_15) begin
      Lsu2Plugin_logic_sq_regs_15_redoSet = 1'b1;
    end
    if(when_Lsu2Plugin_l929) begin
      if(!AguPlugin_setup_port_payload_load) begin
        case(switch_Utils_l1437_3)
          4'b0000 : begin
          end
          4'b0001 : begin
          end
          4'b0010 : begin
          end
          4'b0011 : begin
          end
          4'b0100 : begin
          end
          4'b0101 : begin
          end
          4'b0110 : begin
          end
          4'b0111 : begin
          end
          4'b1000 : begin
          end
          4'b1001 : begin
          end
          4'b1010 : begin
          end
          4'b1011 : begin
          end
          4'b1100 : begin
          end
          4'b1101 : begin
          end
          4'b1110 : begin
          end
          default : begin
            Lsu2Plugin_logic_sq_regs_15_redoSet = 1'b1;
          end
        endcase
      end
    end
    if(Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger) begin
      if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
        if(_zz_134) begin
          Lsu2Plugin_logic_sq_regs_15_redoSet = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_15_delete = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      if(when_Lsu2Plugin_l1524_15) begin
        Lsu2Plugin_logic_sq_regs_15_delete = 1'b1;
      end
    end
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      if(when_Lsu2Plugin_l1909_15) begin
        Lsu2Plugin_logic_sq_regs_15_delete = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_15_commitedNext = Lsu2Plugin_logic_sq_regs_15_commited;
    if(when_Lsu2Plugin_l591) begin
      if(_zz_45[15]) begin
        Lsu2Plugin_logic_sq_regs_15_commitedNext = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l591_1) begin
      if(_zz_46[15]) begin
        Lsu2Plugin_logic_sq_regs_15_commitedNext = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAnySet = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(_zz_134) begin
              Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAnySet = 1'b1;
            end
          end
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign when_Lsu2Plugin_l369_15 = (Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAny && Lsu2Plugin_logic_translationWake);
  assign when_Lsu2Plugin_l385_15 = (Lsu2Plugin_logic_sq_regs_15_redoSet || Lsu2Plugin_logic_sq_regs_15_delete);
  assign Lsu2Plugin_logic_sq_ptr_allocReal = Lsu2Plugin_logic_sq_ptr_alloc[3 : 0];
  assign Lsu2Plugin_logic_sq_ptr_freeReal = Lsu2Plugin_logic_sq_ptr_free[3 : 0];
  assign Lsu2Plugin_logic_sq_ptr_writeBackReal = Lsu2Plugin_logic_sq_ptr_writeBack[3 : 0];
  assign Lsu2Plugin_logic_sq_ptr_commitReal = Lsu2Plugin_logic_sq_ptr_commit[3 : 0];
  assign Lsu2Plugin_logic_sqWritebackEvent_valid = Lsu2Plugin_logic_sq_ptr_onFree_valid;
  assign Lsu2Plugin_logic_sqWritebackEvent_payload = Lsu2Plugin_logic_sq_ptr_onFree_payload;
  assign when_Lsu2Plugin_l572 = (Lsu2Plugin_logic_sq_ptr_commit != Lsu2Plugin_logic_sq_ptr_free);
  assign when_UInt_l120_1 = (|Lsu2Plugin_logic_sq_tracker_freeNext[4 : 2]);
  always @(*) begin
    if(when_UInt_l120_1) begin
      _zz_Lsu2Plugin_logic_sq_tracker_freeReduced = 2'b11;
    end else begin
      _zz_Lsu2Plugin_logic_sq_tracker_freeReduced = Lsu2Plugin_logic_sq_tracker_freeNext[1 : 0];
    end
  end

  assign Lsu2Plugin_logic_sq_tracker_freeNext = (_zz_Lsu2Plugin_logic_sq_tracker_freeNext + _zz_Lsu2Plugin_logic_sq_tracker_freeNext_4);
  assign Lsu2Plugin_logic_sq_onCommit_sqCommits_0 = (CommitPlugin_logic_commit_event_mask[0] && Lsu2Plugin_logic_sq_onCommit_sqAlloc_0);
  assign Lsu2Plugin_logic_sq_onCommit_sqCommits_1 = (CommitPlugin_logic_commit_event_mask[1] && Lsu2Plugin_logic_sq_onCommit_sqAlloc_1);
  assign Lsu2Plugin_logic_sq_onCommit_commitComb = Lsu2Plugin_logic_sq_ptr_commit;
  assign when_Lsu2Plugin_l591 = (CommitPlugin_logic_commit_event_mask[0] && Lsu2Plugin_logic_sq_onCommit_sqAlloc_0);
  assign _zz_45 = ({15'd0,1'b1} <<< Lsu2Plugin_logic_sq_onCommit_commitComb[3 : 0]);
  assign when_Lsu2Plugin_l591_1 = (CommitPlugin_logic_commit_event_mask[1] && Lsu2Plugin_logic_sq_onCommit_sqAlloc_1);
  assign _zz_46 = ({15'd0,1'b1} <<< Lsu2Plugin_logic_sq_onCommit_commitComb_1[3 : 0]);
  assign Lsu2Plugin_logic_sq_ptr_commitNext = Lsu2Plugin_logic_sq_onCommit_commitComb_2;
  always @(*) begin
    FrontendPlugin_dispatch_LSU_ID_0 = 5'bxxxxx;
    if(Lsu2Plugin_logic_allocation_loads_requests_0) begin
      FrontendPlugin_dispatch_LSU_ID_0 = Lsu2Plugin_logic_allocation_loads_alloc;
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_0) begin
      FrontendPlugin_dispatch_LSU_ID_0 = Lsu2Plugin_logic_allocation_stores_alloc;
    end
  end

  always @(*) begin
    FrontendPlugin_dispatch_LSU_ID_1 = 5'bxxxxx;
    if(Lsu2Plugin_logic_allocation_loads_requests_1) begin
      FrontendPlugin_dispatch_LSU_ID_1 = Lsu2Plugin_logic_allocation_loads_alloc_1;
    end
    if(Lsu2Plugin_logic_allocation_stores_requests_1) begin
      FrontendPlugin_dispatch_LSU_ID_1 = Lsu2Plugin_logic_allocation_stores_alloc_1;
    end
  end

  assign Lsu2Plugin_logic_allocation_loads_requests_0 = (FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 && FrontendPlugin_dispatch_LQ_ALLOC_0);
  assign Lsu2Plugin_logic_allocation_loads_requests_1 = (FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1 && FrontendPlugin_dispatch_LQ_ALLOC_1);
  assign Lsu2Plugin_logic_allocation_loads_requestsCount = _zz_Lsu2Plugin_logic_allocation_loads_requestsCount;
  assign Lsu2Plugin_logic_allocation_loads_full = (Lsu2Plugin_logic_lq_tracker_freeReduced < Lsu2Plugin_logic_allocation_loads_requestsCount);
  assign Lsu2Plugin_logic_allocation_loads_alloc = Lsu2Plugin_logic_lq_ptr_alloc;
  assign Lsu2Plugin_logic_allocation_stores_requests_0 = (FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 && FrontendPlugin_dispatch_SQ_ALLOC_0);
  assign Lsu2Plugin_logic_allocation_stores_requests_1 = (FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1 && FrontendPlugin_dispatch_SQ_ALLOC_1);
  assign Lsu2Plugin_logic_allocation_stores_requestsCount = _zz_Lsu2Plugin_logic_allocation_stores_requestsCount;
  assign Lsu2Plugin_logic_allocation_stores_full = (Lsu2Plugin_logic_sq_tracker_freeReduced < Lsu2Plugin_logic_allocation_stores_requestsCount);
  assign Lsu2Plugin_logic_allocation_stores_alloc = Lsu2Plugin_logic_sq_ptr_alloc;
  assign FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l620 = (FrontendPlugin_dispatch_valid && (Lsu2Plugin_logic_allocation_loads_full || Lsu2Plugin_logic_allocation_stores_full));
  assign FrontendPlugin_dispatch_LQ_ID_0 = Lsu2Plugin_logic_allocation_loads_alloc[3:0];
  assign FrontendPlugin_dispatch_SQ_ID_0 = Lsu2Plugin_logic_allocation_stores_alloc[3:0];
  assign FrontendPlugin_dispatch_isFireing = (FrontendPlugin_dispatch_valid && FrontendPlugin_dispatch_ready);
  assign FrontendPlugin_dispatch_LQ_ID_1 = Lsu2Plugin_logic_allocation_loads_alloc_1[3:0];
  assign FrontendPlugin_dispatch_SQ_ID_1 = Lsu2Plugin_logic_allocation_stores_alloc_1[3:0];
  always @(*) begin
    Lsu2Plugin_logic_lq_tracker_sub = 2'b00;
    if(FrontendPlugin_dispatch_isFireing) begin
      Lsu2Plugin_logic_lq_tracker_sub = Lsu2Plugin_logic_allocation_loads_requestsCount;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sq_tracker_sub = 2'b00;
    if(FrontendPlugin_dispatch_isFireing) begin
      Lsu2Plugin_logic_sq_tracker_sub = Lsu2Plugin_logic_allocation_stores_requestsCount;
    end
  end

  assign Lsu2Plugin_logic_aguPush_0_pushLq = (AguPlugin_setup_port_valid && AguPlugin_setup_port_payload_load);
  assign Lsu2Plugin_logic_aguPush_0_pushSq = (AguPlugin_setup_port_valid && (! AguPlugin_setup_port_payload_load));
  always @(*) begin
    _zz_Lsu2Plugin_logic_aguPush_0_dataMask = 4'bxxxx;
    case(AguPlugin_setup_port_payload_size)
      2'b00 : begin
        _zz_Lsu2Plugin_logic_aguPush_0_dataMask = 4'b0001;
      end
      2'b01 : begin
        _zz_Lsu2Plugin_logic_aguPush_0_dataMask = 4'b0011;
      end
      2'b10 : begin
        _zz_Lsu2Plugin_logic_aguPush_0_dataMask = 4'b1111;
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_aguPush_0_dataMask = (_zz_Lsu2Plugin_logic_aguPush_0_dataMask <<< AguPlugin_setup_port_payload_address[1 : 0]);
  assign switch_Utils_l1437 = AguPlugin_setup_port_payload_aguId[3:0];
  assign _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_1 = _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_2;
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score = _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_1[2 : 0];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_tag = _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_1[18 : 3];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_delta = _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_1[22 : 19];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_valid = AguPlugin_setup_port_payload_earlySample;
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_payload = AguPlugin_setup_port_payload_earlyPc[8 : 2];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_hash = AguPlugin_setup_port_payload_pc[24 : 9];
  assign Lsu2Plugin_logic_aguPush_0_hazardPrediction_hit = ((Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score != 3'b000) && (Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_tag == Lsu2Plugin_logic_aguPush_0_hazardPrediction_hash));
  assign Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter = _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter_1[5 : 0];
  assign Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_valid = AguPlugin_setup_port_payload_earlySample;
  assign Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_payload = AguPlugin_setup_port_payload_earlyPc[11 : 2];
  assign Lsu2Plugin_logic_aguPush_0_hitPrediction_likelyToHit = Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter[5];
  assign when_Lsu2Plugin_l733 = (Lsu2Plugin_logic_aguPush_0_pushSq && (AguPlugin_setup_port_payload_sc || AguPlugin_setup_port_payload_amo));
  assign switch_Utils_l1437_1 = AguPlugin_setup_port_payload_aguId[3:0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo = {Lsu2Plugin_logic_lq_regs_15_redo,{Lsu2Plugin_logic_lq_regs_14_redo,{Lsu2Plugin_logic_lq_regs_13_redo,{Lsu2Plugin_logic_lq_regs_12_redo,{Lsu2Plugin_logic_lq_regs_11_redo,{Lsu2Plugin_logic_lq_regs_10_redo,{Lsu2Plugin_logic_lq_regs_9_redo,{Lsu2Plugin_logic_lq_regs_8_redo,{Lsu2Plugin_logic_lq_regs_7_redo,{Lsu2Plugin_logic_lq_regs_6_redo,{_zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo,_zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_1}}}}}}}}}}};
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo = {Lsu2Plugin_logic_sq_regs_15_redo,{Lsu2Plugin_logic_sq_regs_14_redo,{Lsu2Plugin_logic_sq_regs_13_redo,{Lsu2Plugin_logic_sq_regs_12_redo,{Lsu2Plugin_logic_sq_regs_11_redo,{Lsu2Plugin_logic_sq_regs_10_redo,{Lsu2Plugin_logic_sq_regs_9_redo,{Lsu2Plugin_logic_sq_regs_8_redo,{Lsu2Plugin_logic_sq_regs_7_redo,{Lsu2Plugin_logic_sq_regs_6_redo,{_zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo,_zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_1}}}}}}}}}}};
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_input = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_priorityBits = Lsu2Plugin_logic_lq_ptr_priority;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask = {Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_input,(Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_input[15 : 1] & Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_priorityBits)};
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0 = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_1 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[1];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_2 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[2];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[3];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[4];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_5 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[5];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[6];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_7 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[7];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_8 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[8];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[9];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[10];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_11 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[11];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[12];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_13 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[13];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_14 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[14];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_15 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[15];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_16 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[16];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_17 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[17];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_18 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[18];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_19 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[19];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_20 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[20];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_21 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[21];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_22 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[22];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_23 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[23];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_24 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[24];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_25 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[25];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_26 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[26];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_27 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[27];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_28 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[28];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_29 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[29];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_30 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0[30];
  always @(*) begin
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[0] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[1] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_1 && (! Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[2] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_2 && (! Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[3] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3 && (! Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[4] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[5] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_5 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_4 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[6] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_5 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[7] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_7 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[8] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_8 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_7 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[9] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_8 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[10] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[11] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_11 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_9_to_10 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[12] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_9_to_11 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[13] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_13 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[14] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_14 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_13 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[15] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_15 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_14 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[16] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_16 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_15 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[17] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_17 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_15_to_16 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[18] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_18 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_15_to_17 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[19] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_19 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_18 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[20] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_20 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_19 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[21] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_21 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[22] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_22 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_21 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[23] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_23 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_21_to_22 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[24] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_24 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_21_to_23 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[25] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_25 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_24 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[26] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_26 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_24_to_25 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[27] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_27 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_24_to_26 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[28] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_28 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_27 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[29] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_29 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_27_to_28 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[30] = (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_30 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_27_to_29 || (Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
  end

  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_1 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_2,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_0}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_4 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_5 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_5,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_4,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_3}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_5 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_7 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_8 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_8,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_6}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_8 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_9_to_10 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_9_to_11 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_11,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_10,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_9}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_11 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2}}} != 4'b0000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_13 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_14 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_14,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_12}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_14 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_14,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2}}}} != 5'h00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_15_to_16 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_16,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_15} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_15_to_17 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_17,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_16,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_15}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_17 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_15_to_17,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_12_to_14,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_0_to_2}}}}} != 6'h00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_19 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_19,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_18} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_20 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_20,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_19,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_18}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_21_to_22 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_22,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_21} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_21_to_23 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_23,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_22,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_21}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_23 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_21_to_23,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_20} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_24_to_25 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_25,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_24} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_24_to_26 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_26,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_25,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_24}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_26 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_24_to_26,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_21_to_23,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_18_to_20}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_27_to_28 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_28,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_27} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_range_27_to_29 = ({Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_29,{Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_28,Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleMask_bools_27}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pLow = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[30 : 15];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pHigh = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_doubleOh[14 : 0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh = (_zz_Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh | Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_pLow);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH = Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo_roundRobinMasked_selOh;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_input = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_priorityBits = Lsu2Plugin_logic_sq_ptr_priority;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask = {Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_input,(Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_input[15 : 1] & Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_priorityBits)};
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0 = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_1 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[1];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_2 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[2];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[3];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[4];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_5 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[5];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[6];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_7 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[7];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_8 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[8];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[9];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[10];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_11 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[11];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[12];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_13 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[13];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_14 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[14];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_15 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[15];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_16 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[16];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_17 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[17];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_18 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[18];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_19 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[19];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_20 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[20];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_21 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[21];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_22 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[22];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_23 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[23];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_24 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[24];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_25 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[25];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_26 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[26];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_27 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[27];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_28 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[28];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_29 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[29];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_30 = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0[30];
  always @(*) begin
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[0] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[1] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_1 && (! Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[2] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_2 && (! Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[3] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3 && (! Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[4] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[5] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_5 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_4 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[6] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_5 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[7] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_7 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[8] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_8 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_7 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[9] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_8 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[10] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[11] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_11 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_9_to_10 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[12] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_9_to_11 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[13] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_13 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[14] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_14 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_13 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[15] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_15 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_14 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[16] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_16 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_15 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[17] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_17 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_15_to_16 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[18] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_18 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_15_to_17 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[19] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_19 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_18 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[20] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_20 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_19 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[21] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_21 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[22] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_22 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_21 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[23] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_23 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_21_to_22 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[24] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_24 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_21_to_23 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[25] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_25 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_24 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[26] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_26 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_24_to_25 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[27] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_27 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_24_to_26 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[28] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_28 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_27 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[29] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_29 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_27_to_28 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[30] = (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_30 && (! (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_27_to_29 || (Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17))));
  end

  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_1 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_2,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_0}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_4 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_5 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_5,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_4,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_3}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_5 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_7 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_8 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_8,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_6}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_8 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_9_to_10 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_9_to_11 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_11,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_10,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_9}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_11 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2}}} != 4'b0000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_13 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_14 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_14,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_12}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_14 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_14,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2}}}} != 5'h00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_15_to_16 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_16,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_15} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_15_to_17 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_17,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_16,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_15}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_17 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_15_to_17,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_12_to_14,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_0_to_2}}}}} != 6'h00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_19 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_19,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_18} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_20 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_20,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_19,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_18}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_21_to_22 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_22,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_21} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_21_to_23 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_23,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_22,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_21}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_23 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_21_to_23,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_20} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_24_to_25 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_25,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_24} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_24_to_26 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_26,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_25,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_24}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_26 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_24_to_26,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_21_to_23,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_18_to_20}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_27_to_28 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_28,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_27} != 2'b00);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_range_27_to_29 = ({Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_29,{Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_28,Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleMask_bools_27}} != 3'b000);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh = _zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pLow = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[30 : 15];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pHigh = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_doubleOh[14 : 0];
  assign Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh = (_zz_Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh | Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_pLow);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH = Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo_roundRobinMasked_selOh;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT = (|Lsu2Plugin_logic_lqSqArbitration_s0_lqRedo);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT = (|Lsu2Plugin_logic_lqSqArbitration_s0_sqRedo);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[1];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_1 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[2];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[3];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_3 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[4];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[5];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[6];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[7];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_7 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[8];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_8 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[9];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_9 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[10];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_10 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[11];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_11 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[12];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_12 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[13];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_13 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[14];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_14 = Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[15];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_15 = (((((((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_8) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_10) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_12) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_14);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_16 = (((((((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_1 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_9) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_10) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_13) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_14);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_17 = (((((((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_3 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_11) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_12) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_13) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_14);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_18 = (((((((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_7 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_8) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_9) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_10) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_11) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_12) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_13) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_14);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID = {_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_18,{_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_17,{_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_16,_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_15}}};
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[1];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_1 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[2];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[3];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_3 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[4];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[5];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[6];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[7];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_7 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[8];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_8 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[9];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_9 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[10];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_10 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[11];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_11 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[12];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_12 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[13];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_13 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[14];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_14 = Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[15];
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_15 = (((((((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_8) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_10) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_12) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_14);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_16 = (((((((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_1 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_9) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_10) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_13) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_14);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_17 = (((((((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_3 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_11) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_12) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_13) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_14);
  assign _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_18 = (((((((_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_7 || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_8) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_9) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_10) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_11) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_12) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_13) || _zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_14);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID = {_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_18,{_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_17,{_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_16,_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_15}}};
  assign Lsu2Plugin_logic_lqSqArbitration_s0_valid = (Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT || Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT);
  assign Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ROB_FULL = {_zz_Lsu2Plugin_logic_lq_mem_robIdMsb_port1,_zz_Lsu2Plugin_logic_lq_mem_robId_port1};
  assign Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ROB_FULL = {_zz_Lsu2Plugin_logic_sq_mem_robIdMsb_port1,_zz_Lsu2Plugin_logic_sq_mem_robId_port1};
  assign Lsu2Plugin_logic_lqSqArbitration_s1_cmp = _zz_Lsu2Plugin_logic_lqSqArbitration_s1_cmp[6];
  assign Lsu2Plugin_logic_lqSqArbitration_s1_LQ_OLDER_THAN_SQ = ((! Lsu2Plugin_logic_lqSqArbitration_s1_SQ_HIT) || (Lsu2Plugin_logic_lqSqArbitration_s1_LQ_HIT && Lsu2Plugin_logic_lqSqArbitration_s1_cmp));
  assign Lsu2Plugin_logic_translationWake = Lsu2Plugin_logic_sharedPip_translationPort_wake;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION) begin
        Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_speculateHitTrapRecovered = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            Lsu2Plugin_logic_sharedPip_speculateHitTrapRecovered = (Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID == 4'b0000);
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION = 1'b0;
    if(when_Lsu2Plugin_l920) begin
      Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ = Lsu2Plugin_logic_lqSqArbitration_s1_LQ_OLDER_THAN_SQ;
    if(when_Lsu2Plugin_l838) begin
      Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ = 1'b0;
    end
    if(when_Lsu2Plugin_l839) begin
      Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_LQ_ROB_FULL = Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ROB_FULL;
  assign Lsu2Plugin_logic_sharedPip_stages_0_SQ_ROB_FULL = Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ROB_FULL;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_feed_takeAgu = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu[6] : _zz_Lsu2Plugin_logic_sharedPip_feed_takeAgu_1[6]);
    if(when_Lsu2Plugin_l830) begin
      Lsu2Plugin_logic_sharedPip_feed_takeAgu = 1'b1;
    end
    if(when_Lsu2Plugin_l831) begin
      Lsu2Plugin_logic_sharedPip_feed_takeAgu = 1'b0;
    end
  end

  assign when_Lsu2Plugin_l830 = (! Lsu2Plugin_logic_lqSqArbitration_s1_valid);
  assign when_Lsu2Plugin_l831 = (! AguPlugin_setup_port_valid);
  assign Lsu2Plugin_logic_sharedPip_stages_0_valid = (AguPlugin_setup_port_valid || Lsu2Plugin_logic_lqSqArbitration_s1_valid);
  assign Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l834 = (Lsu2Plugin_logic_sharedPip_feed_takeAgu || (! Lsu2Plugin_logic_sharedPip_stages_0_ready));
  assign when_Lsu2Plugin_l838 = (! Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask);
  assign when_Lsu2Plugin_l839 = (! Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask);
  assign when_Lsu2Plugin_l841 = (((Lsu2Plugin_logic_lqSqArbitration_s1_SQ_HIT && Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask) && Lsu2Plugin_logic_lqSqArbitration_s1_LQ_HIT) && Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask);
  assign Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842 = _zz_Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842;
  assign when_Lsu2Plugin_l843 = ((! Lsu2Plugin_logic_sharedPip_feed_takeAgu) && Lsu2Plugin_logic_sharedPip_stages_0_ready);
  assign when_Lsu2Plugin_l845 = (! Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ);
  assign when_Lsu2Plugin_l849 = ((Lsu2Plugin_logic_lqSqArbitration_s1_isRemoved || Lsu2Plugin_logic_lqSqArbitration_s1_ready) || (! Lsu2Plugin_logic_lqSqArbitration_s1_valid));
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID = _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID[5:0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID = _zz_Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_1[5:0];
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD = _zz_Lsu2Plugin_logic_lq_mem_physRd_port1;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD = AguPlugin_setup_port_payload_physicalRd;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_load = _zz_Lsu2Plugin_logic_lq_mem_addressPre_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_store = _zz_Lsu2Plugin_logic_sq_mem_addressPre_port1;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_load : Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION_store);
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION = AguPlugin_setup_port_payload_address;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_load = _zz_Lsu2Plugin_logic_lq_mem_addressPost_port0;
  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_store = _zz_Lsu2Plugin_logic_sq_mem_addressPost_port0;
  assign Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_load : Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION_store);
  assign Lsu2Plugin_logic_sharedPip_stages_0_SIZE_load = _zz_Lsu2Plugin_logic_lq_mem_size_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_SIZE_store = _zz_Lsu2Plugin_logic_sq_mem_size_port1;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_SIZE = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_SIZE_load : Lsu2Plugin_logic_sharedPip_stages_0_SIZE_store);
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_SIZE = AguPlugin_setup_port_payload_size;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_load = Lsu2Plugin_logic_lq_mem_needTranslation_io_read_0_rsp[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_store = Lsu2Plugin_logic_sq_mem_needTranslation_io_read_0_rsp[0];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_load : Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION_store);
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_load = _zz_Lsu2Plugin_logic_lq_mem_io_port0[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_store = _zz_Lsu2Plugin_logic_sq_mem_io_port0[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO = (Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ ? Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_load : Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO_store);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD = _zz_Lsu2Plugin_logic_lq_mem_writeRd_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD = AguPlugin_setup_port_payload_writeRd;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_UNSIGNED = _zz_Lsu2Plugin_logic_lq_mem_unsigned_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_UNSIGNED = AguPlugin_setup_port_payload_unsigned;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LR = _zz_Lsu2Plugin_logic_lq_mem_lr_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LR = AguPlugin_setup_port_payload_lr;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC = Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_0_rsp;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LQ_SQ_ALLOC = Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_1_rsp;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID = _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_valid_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID = Lsu2Plugin_logic_aguPush_0_hazardPrediction_hit;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA = _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_delta_port1;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA = Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_delta;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SCORE = _zz_Lsu2Plugin_logic_lq_mem_hazardPrediction_score_port1;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SCORE = Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_AMO = _zz_Lsu2Plugin_logic_sq_mem_amo_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_AMO = AguPlugin_setup_port_payload_amo;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_SC = _zz_Lsu2Plugin_logic_sq_mem_sc_port1[0];
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_SC = AguPlugin_setup_port_payload_sc;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD = Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD = AguPlugin_setup_port_payload_load;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID = Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID = AguPlugin_setup_port_payload_aguId[3:0];
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID = Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID = AguPlugin_setup_port_payload_aguId[3:0];
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_feed_takeAgu) begin
      Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION_COUNTER = Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter;
  assign Lsu2Plugin_logic_sharedPip_stages_0_SP_FP_ADDRESS = 1'b0;
  assign when_Lsu2Plugin_l920 = ((((! Lsu2Plugin_logic_lqSqArbitration_s1_valid) && AguPlugin_setup_port_payload_load) && (Lsu2Plugin_logic_aguPush_0_hitPrediction_likelyToHit || Lsu2Plugin_logic_sharedPip_stages_0_SP_FP_ADDRESS)) && Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled);
  assign Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_agu = AguPlugin_setup_port_payload_robId;
  assign Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD_agu = AguPlugin_setup_port_payload_writeRd;
  assign Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD_agu = AguPlugin_setup_port_payload_physicalRd;
  assign when_Lsu2Plugin_l929 = (AguPlugin_setup_port_valid && ((! Lsu2Plugin_logic_sharedPip_feed_takeAgu) || (! Lsu2Plugin_logic_sharedPip_stages_0_ready)));
  assign switch_Utils_l1437_2 = AguPlugin_setup_port_payload_aguId[3:0];
  assign switch_Utils_l1437_3 = AguPlugin_setup_port_payload_aguId[3:0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_isFireing = (Lsu2Plugin_logic_sharedPip_stages_0_valid && Lsu2Plugin_logic_sharedPip_stages_0_ready);
  assign Lsu2Plugin_logic_sqFeedEvent_valid = (Lsu2Plugin_logic_sharedPip_stages_0_isFireing && (! Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD));
  assign Lsu2Plugin_logic_sqFeedEvent_payload = Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID;
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = 4'bxxxx;
    case(Lsu2Plugin_logic_sharedPip_stages_0_SIZE)
      2'b00 : begin
        _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = 4'b0001;
      end
      2'b01 : begin
        _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = 4'b0011;
      end
      2'b10 : begin
        _zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = 4'b1111;
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK = (_zz_Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK <<< Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[1 : 0]);
  assign Lsu2Plugin_logic_sharedPip_stages_0_LQCHECK_START_ID = Lsu2Plugin_logic_sq_mem_lqAlloc_io_read_0_rsp;
  assign Lsu2Plugin_logic_sharedPip_stages_0_SQCHECK_END_ID = Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_2_rsp;
  assign Lsu2Plugin_logic_sharedPip_stages_0_feed_SQ_PTR_FREE = Lsu2Plugin_logic_sq_ptr_free;
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT = (_zz__zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT - 5'h01);
  assign Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SQID = _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT[3:0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT = ((Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID && (! Lsu2Plugin_logic_sq_mem_feededOnce_io_read_0_rsp[0])) && (! _zz_Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_1[4]));
  assign Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_FEEDED = 1'b0;
  assign Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded = (Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED || (Lsu2Plugin_logic_sqFeedEvent_valid && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SQID)));
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded = (Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED || (Lsu2Plugin_logic_sqFeedEvent_valid && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SQID)));
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED || (Lsu2Plugin_logic_sqFeedEvent_valid && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SQID)));
  assign Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH_PC = AguPlugin_setup_port_payload_pc;
  assign when_Lsu2Plugin_l959 = (Lsu2Plugin_logic_sharedPip_stages_0_isFireing && (! Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD));
  assign Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_valid = (Lsu2Plugin_logic_sharedPip_stages_0_isFireing && Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION);
  assign Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_payload_robId = Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID_agu;
  assign Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_valid = ((Lsu2Plugin_logic_sharedPip_stages_0_isFireing && Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION) && Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD_agu);
  assign Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_payload_physical = Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD_agu;
  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_valid = (Lsu2Plugin_logic_sharedPip_stages_0_valid != 1'b0);
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_valid = 1'b1;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_payload_virtual = Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_payload_virtual = Lsu2Plugin_logic_special_storeAddress;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_payload_size = Lsu2Plugin_logic_sharedPip_stages_0_SIZE;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_payload_size = Lsu2Plugin_logic_special_storeSize;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_payload_redoOnDataHazard = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_payload_redoOnDataHazard = 1'b0;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_cmd_payload_unique = ((! Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD) || Lsu2Plugin_logic_sharedPip_stages_0_LR);
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
        Lsu2Plugin_setup_cacheLoad_cmd_payload_unique = 1'b1;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_haltRequest_Lsu2Plugin_l990 = (! Lsu2Plugin_setup_cacheLoad_cmd_ready);
  assign when_Lsu2Plugin_l997 = (! Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION);
  always @(*) begin
    if(when_Lsu2Plugin_l997) begin
      Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_POST_TRANSLATION;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED = Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
    end
  end

  always @(*) begin
    if(when_Lsu2Plugin_l997) begin
      Lsu2Plugin_logic_sharedPip_stages_1_IS_IO = Lsu2Plugin_logic_sharedPip_stages_1_TRANSLATED_AS_IO;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_IS_IO = Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_translated_physical = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED;
    if(when_Lsu2Plugin_l1683) begin
      Lsu2Plugin_setup_cacheLoad_translated_physical = Lsu2Plugin_logic_special_storeAddress;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheLoad_translated_abord = (Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION ? ((((Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO || Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT) || Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT) || (! Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ)) || Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO) : Lsu2Plugin_logic_sharedPip_stages_1_TRANSLATED_AS_IO);
    if(when_Lsu2Plugin_l1683) begin
      Lsu2Plugin_setup_cacheLoad_translated_abord = 1'b0;
    end
  end

  assign Lsu2Plugin_setup_cacheLoad_cancels = 3'b000;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask = Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE[3 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask = {1'b0,{(4'b1110 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(4'b1101 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(4'b1100 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(4'b1011 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_1 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask),{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_2,{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_3,_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask_4}}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID[3 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask = {1'b0,{(4'b1110 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(4'b1101 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(4'b1100 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(4'b1011 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_1 < _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask),{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_2,{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_3,_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask_4}}}}}}}};
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_loopback = (Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE[4] != Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID[4]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_youngerMask = (Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_loopback ? (~ (Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask ^ Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask)) : (Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_endMask & (~ Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_startMask)));
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_olderMaskEmpty = (Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE == Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK = Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_youngerMask;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_NO_OLDER = Lsu2Plugin_logic_sharedPip_checkSqMask_maskGen_olderMaskEmpty;
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_pageHit = (Lsu2Plugin_logic_sq_regs_0_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_wordHit = ((Lsu2Plugin_logic_sq_regs_0_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[0] = ((((Lsu2Plugin_logic_sq_regs_0_valid && Lsu2Plugin_logic_sq_regs_0_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_0_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[0]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[1] = ((((Lsu2Plugin_logic_sq_regs_1_valid && Lsu2Plugin_logic_sq_regs_1_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[1]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[2] = ((((Lsu2Plugin_logic_sq_regs_2_valid && Lsu2Plugin_logic_sq_regs_2_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[2]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[3] = ((((Lsu2Plugin_logic_sq_regs_3_valid && Lsu2Plugin_logic_sq_regs_3_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[3]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[4] = ((((Lsu2Plugin_logic_sq_regs_4_valid && Lsu2Plugin_logic_sq_regs_4_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[4]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[5] = ((((Lsu2Plugin_logic_sq_regs_5_valid && Lsu2Plugin_logic_sq_regs_5_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[5]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[6] = ((((Lsu2Plugin_logic_sq_regs_6_valid && Lsu2Plugin_logic_sq_regs_6_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[6]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[7] = ((((Lsu2Plugin_logic_sq_regs_7_valid && Lsu2Plugin_logic_sq_regs_7_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[7]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[8] = ((((Lsu2Plugin_logic_sq_regs_8_valid && Lsu2Plugin_logic_sq_regs_8_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_8_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_8_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[8]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[9] = ((((Lsu2Plugin_logic_sq_regs_9_valid && Lsu2Plugin_logic_sq_regs_9_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_9_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_9_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[9]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[10] = ((((Lsu2Plugin_logic_sq_regs_10_valid && Lsu2Plugin_logic_sq_regs_10_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_10_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_10_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[10]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[11] = ((((Lsu2Plugin_logic_sq_regs_11_valid && Lsu2Plugin_logic_sq_regs_11_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_11_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_11_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[11]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[12] = ((((Lsu2Plugin_logic_sq_regs_12_valid && Lsu2Plugin_logic_sq_regs_12_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_12_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_12_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[12]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[13] = ((((Lsu2Plugin_logic_sq_regs_13_valid && Lsu2Plugin_logic_sq_regs_13_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_13_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_13_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[13]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[14] = ((((Lsu2Plugin_logic_sq_regs_14_valid && Lsu2Plugin_logic_sq_regs_14_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_14_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_14_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[14]);
    Lsu2Plugin_logic_sharedPip_checkSqMask_hits[15] = ((((Lsu2Plugin_logic_sq_regs_15_valid && Lsu2Plugin_logic_sq_regs_15_dataValid) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_15_pageHit) && Lsu2Plugin_logic_sharedPip_checkSqMask_entries_15_wordHit) && Lsu2Plugin_logic_sharedPip_stages_1_SQ_YOUNGER_MASK[15]);
  end

  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_pageHit = (Lsu2Plugin_logic_sq_regs_1_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_1_wordHit = ((Lsu2Plugin_logic_sq_regs_1_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_pageHit = (Lsu2Plugin_logic_sq_regs_2_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_2_wordHit = ((Lsu2Plugin_logic_sq_regs_2_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_pageHit = (Lsu2Plugin_logic_sq_regs_3_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_3_wordHit = ((Lsu2Plugin_logic_sq_regs_3_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_pageHit = (Lsu2Plugin_logic_sq_regs_4_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_4_wordHit = ((Lsu2Plugin_logic_sq_regs_4_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_pageHit = (Lsu2Plugin_logic_sq_regs_5_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_5_wordHit = ((Lsu2Plugin_logic_sq_regs_5_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_pageHit = (Lsu2Plugin_logic_sq_regs_6_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_6_wordHit = ((Lsu2Plugin_logic_sq_regs_6_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_pageHit = (Lsu2Plugin_logic_sq_regs_7_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_7_wordHit = ((Lsu2Plugin_logic_sq_regs_7_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_8_pageHit = (Lsu2Plugin_logic_sq_regs_8_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_8_wordHit = ((Lsu2Plugin_logic_sq_regs_8_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_9_pageHit = (Lsu2Plugin_logic_sq_regs_9_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_9_wordHit = ((Lsu2Plugin_logic_sq_regs_9_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_10_pageHit = (Lsu2Plugin_logic_sq_regs_10_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_10_wordHit = ((Lsu2Plugin_logic_sq_regs_10_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_11_pageHit = (Lsu2Plugin_logic_sq_regs_11_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_11_wordHit = ((Lsu2Plugin_logic_sq_regs_11_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_12_pageHit = (Lsu2Plugin_logic_sq_regs_12_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_12_wordHit = ((Lsu2Plugin_logic_sq_regs_12_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_13_pageHit = (Lsu2Plugin_logic_sq_regs_13_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_13_wordHit = ((Lsu2Plugin_logic_sq_regs_13_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_14_pageHit = (Lsu2Plugin_logic_sq_regs_14_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_14_wordHit = ((Lsu2Plugin_logic_sq_regs_14_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_15_pageHit = (Lsu2Plugin_logic_sq_regs_15_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_entries_15_wordHit = ((Lsu2Plugin_logic_sq_regs_15_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS = Lsu2Plugin_logic_sharedPip_checkSqMask_hits;
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_olderHit = ((! Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_NO_OLDER) && (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS != 16'h0000));
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input = {_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[0],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[1],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[2],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[3],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[4],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[5],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[6],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input_1,{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input_2,_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input_3}}}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits = Lsu2Plugin_logic_sq_ptr_priorityLast;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits = (~ {_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[0],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[1],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[2],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[3],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[4],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[5],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits[6],{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits_1,{_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits_2,_zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits_3}}}}}}}}});
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask = {{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[14 : 0],Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[15 : 15]},(Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_input[14 : 0] & Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_priorityBits)};
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[0];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_1 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[1];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[2];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[3];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[4];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_5 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[5];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[6];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_7 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[7];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[8];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[9];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[10];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_11 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[11];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[12];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_13 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[13];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_14 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[14];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_15 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[15];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_16 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[16];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_17 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[17];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_18 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[18];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_19 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[19];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_20 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[20];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_21 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[21];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_22 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[22];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_23 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[23];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_24 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[24];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_25 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[25];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_26 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[26];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_27 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[27];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_28 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[28];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_29 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[29];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_30 = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[30];
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[0] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[1] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_1 && (! Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[2] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 && (! Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[3] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 && (! Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[4] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[5] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_5 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_4 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[6] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[7] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_7 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[8] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[9] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[10] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[11] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_11 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_10 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[12] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[13] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_13 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[14] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_14 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[15] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_15 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[16] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_16 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_15 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[17] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_17 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_16 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[18] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_18 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_17 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[19] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_19 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_18 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[20] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_20 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_19 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[21] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_21 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[22] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_22 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_21 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[23] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_23 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_22 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[24] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_24 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[25] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_25 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_24 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[26] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_26 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_25 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[27] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_27 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_26 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[28] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_28 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_27 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[29] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_29 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_28 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[30] = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_30 && (! (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_29 || (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
  end

  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_2,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_0}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_4 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_5,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_4,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_3}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_8,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_6}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_10 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_11,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_10,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_9}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2}}} != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_14,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_12}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2}}}} != 5'h00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_16 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_16,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_15} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_17 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_17,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_16,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_15}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_17,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2}}}}} != 6'h00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_19 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_19,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_18} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_20,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_19,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_18}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_22 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_22,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_21} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_23,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_22,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_21}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_25 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_25,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_24} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_26 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_26,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_25,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_24}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_26,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_28 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_28,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_27} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_29 = ({Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_29,{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_28,Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleMask_bools_27}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh = _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh;
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pLow = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[30 : 16];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pHigh = Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_doubleOh[15 : 0];
  assign Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh = (Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_pHigh | _zz_Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh = {Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[0],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[1],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[2],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[3],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[4],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[5],{Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_HITS_roundRobinMasked_selOh[6],{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh,{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh_1,_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh_2}}}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[3];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_1 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[5];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_2 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[6];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[7];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_4 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[9];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_5 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[10];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_6 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[11];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_7 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[12];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_8 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[13];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_9 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[14];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_10 = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[15];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_11 = (((((((Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[1] || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_1) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_4) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_6) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_8) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_10);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_12 = (((((((Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[2] || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_2) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_5) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_6) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_9) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_10);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_13 = (((((((Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[4] || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_1) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_2) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_3) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_7) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_8) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_9) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_10);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_14 = (((((((Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh[8] || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_4) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_5) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_6) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_7) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_8) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_9) || _zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_10);
  assign Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel = {_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_14,{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_13,{_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_12,_zz_Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel_11}}};
  assign Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_HIT = Lsu2Plugin_logic_sharedPip_checkSqMask_olderHit;
  assign Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_ID = Lsu2Plugin_logic_sharedPip_checkSqMask_olderSel;
  assign Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_OH = Lsu2Plugin_logic_sharedPip_checkSqMask_olderOh;
  assign Lsu2Plugin_logic_sharedPip_stages_1_isFireing = (Lsu2Plugin_logic_sharedPip_stages_1_valid && Lsu2Plugin_logic_sharedPip_stages_1_ready);
  assign when_Lsu2Plugin_l1046 = ((Lsu2Plugin_logic_sharedPip_stages_1_isFireing && Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD) && (! Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT));
  assign when_Lsu2Plugin_l1052 = (Lsu2Plugin_logic_sharedPip_stages_1_isFireing && Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION);
  assign Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED = (Lsu2Plugin_logic_sq_ptr_onFreeLast_valid && (Lsu2Plugin_logic_sq_ptr_onFreeLast_payload == Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID));
  assign Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED_overloaded = ((Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED || (Lsu2Plugin_logic_sq_ptr_onFree_valid && (Lsu2Plugin_logic_sq_ptr_onFree_payload == Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID))) || ((Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID)));
  assign Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_overloaded = ((Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED || (Lsu2Plugin_logic_sq_ptr_onFree_valid && (Lsu2Plugin_logic_sq_ptr_onFree_payload == Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID))) || ((Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED && Lsu2Plugin_logic_sqFeedEvent_valid) && (Lsu2Plugin_logic_sqFeedEvent_payload == Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID)));
  assign Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_addressMatch = (_zz_Lsu2Plugin_logic_sq_mem_addressPost_port2 == Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_TRANSLATED);
  assign Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_fullMatch = ((Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_addressMatch && (_zz_Lsu2Plugin_logic_sq_mem_size_port2 == Lsu2Plugin_logic_sharedPip_stages_2_SIZE)) && (! _zz_Lsu2Plugin_logic_sq_mem_doNotBypass_port1[0]));
  assign Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_translationFailure = Lsu2Plugin_logic_sq_mem_needTranslation_io_read_1_rsp[0];
  assign Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_data = _zz_Lsu2Plugin_logic_sq_mem_data_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_BYPASS_SUCCESS = ((! Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_translationFailure) && Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_fullMatch);
  assign Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED = Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_translationFailure;
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_endId = Lsu2Plugin_logic_lq_ptr_alloc;
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask = Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID[3 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_startMask = {1'b0,{(4'b1110 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(4'b1101 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(4'b1100 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(4'b1011 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_1 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask),{_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_2,{_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_3,_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_startMask_4}}}}}}}};
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask = Lsu2Plugin_logic_sharedPip_checkLqHits_endId[3 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_endMask = {1'b0,{(4'b1110 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(4'b1101 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(4'b1100 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(4'b1011 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{(_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_1 < _zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask),{_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_2,{_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_3,_zz_Lsu2Plugin_logic_sharedPip_checkLqHits_endMask_4}}}}}}}};
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_loopback = (Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID[4] != Lsu2Plugin_logic_sharedPip_checkLqHits_endId[4]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask = (Lsu2Plugin_logic_sharedPip_checkLqHits_loopback ? (~ (Lsu2Plugin_logic_sharedPip_checkLqHits_endMask ^ Lsu2Plugin_logic_sharedPip_checkLqHits_startMask)) : (Lsu2Plugin_logic_sharedPip_checkLqHits_endMask & (~ Lsu2Plugin_logic_sharedPip_checkLqHits_startMask)));
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMaskEmpty = (Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID == Lsu2Plugin_logic_sharedPip_checkLqHits_endId);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_pageHit = (Lsu2Plugin_logic_lq_regs_0_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_wordHit = ((Lsu2Plugin_logic_lq_regs_0_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_hit = ((((Lsu2Plugin_logic_lq_regs_0_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_wordHit) && Lsu2Plugin_logic_lq_regs_0_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[0]);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[0] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_hit && Lsu2Plugin_logic_lq_regs_0_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[1] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_hit && Lsu2Plugin_logic_lq_regs_1_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[2] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_hit && Lsu2Plugin_logic_lq_regs_2_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[3] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_hit && Lsu2Plugin_logic_lq_regs_3_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[4] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_hit && Lsu2Plugin_logic_lq_regs_4_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[5] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_hit && Lsu2Plugin_logic_lq_regs_5_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[6] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_hit && Lsu2Plugin_logic_lq_regs_6_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[7] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_hit && Lsu2Plugin_logic_lq_regs_7_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[8] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_hit && Lsu2Plugin_logic_lq_regs_8_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[9] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_hit && Lsu2Plugin_logic_lq_regs_9_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[10] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_hit && Lsu2Plugin_logic_lq_regs_10_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[11] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_hit && Lsu2Plugin_logic_lq_regs_11_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[12] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_hit && Lsu2Plugin_logic_lq_regs_12_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[13] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_hit && Lsu2Plugin_logic_lq_regs_13_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[14] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_hit && Lsu2Plugin_logic_lq_regs_14_sqChecked);
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS[15] = (Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_hit && Lsu2Plugin_logic_lq_regs_15_sqChecked);
  end

  assign when_Lsu2Plugin_l1104 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_0_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_pageHit = (Lsu2Plugin_logic_lq_regs_1_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_wordHit = ((Lsu2Plugin_logic_lq_regs_1_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_hit = ((((Lsu2Plugin_logic_lq_regs_1_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_wordHit) && Lsu2Plugin_logic_lq_regs_1_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[1]);
  assign when_Lsu2Plugin_l1104_1 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_1_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_pageHit = (Lsu2Plugin_logic_lq_regs_2_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_wordHit = ((Lsu2Plugin_logic_lq_regs_2_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_hit = ((((Lsu2Plugin_logic_lq_regs_2_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_wordHit) && Lsu2Plugin_logic_lq_regs_2_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[2]);
  assign when_Lsu2Plugin_l1104_2 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_2_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_pageHit = (Lsu2Plugin_logic_lq_regs_3_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_wordHit = ((Lsu2Plugin_logic_lq_regs_3_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_hit = ((((Lsu2Plugin_logic_lq_regs_3_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_wordHit) && Lsu2Plugin_logic_lq_regs_3_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[3]);
  assign when_Lsu2Plugin_l1104_3 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_3_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_pageHit = (Lsu2Plugin_logic_lq_regs_4_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_wordHit = ((Lsu2Plugin_logic_lq_regs_4_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_hit = ((((Lsu2Plugin_logic_lq_regs_4_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_wordHit) && Lsu2Plugin_logic_lq_regs_4_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[4]);
  assign when_Lsu2Plugin_l1104_4 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_4_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_pageHit = (Lsu2Plugin_logic_lq_regs_5_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_wordHit = ((Lsu2Plugin_logic_lq_regs_5_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_hit = ((((Lsu2Plugin_logic_lq_regs_5_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_wordHit) && Lsu2Plugin_logic_lq_regs_5_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[5]);
  assign when_Lsu2Plugin_l1104_5 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_5_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_pageHit = (Lsu2Plugin_logic_lq_regs_6_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_wordHit = ((Lsu2Plugin_logic_lq_regs_6_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_hit = ((((Lsu2Plugin_logic_lq_regs_6_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_wordHit) && Lsu2Plugin_logic_lq_regs_6_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[6]);
  assign when_Lsu2Plugin_l1104_6 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_6_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_pageHit = (Lsu2Plugin_logic_lq_regs_7_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_wordHit = ((Lsu2Plugin_logic_lq_regs_7_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_hit = ((((Lsu2Plugin_logic_lq_regs_7_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_wordHit) && Lsu2Plugin_logic_lq_regs_7_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[7]);
  assign when_Lsu2Plugin_l1104_7 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_7_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_pageHit = (Lsu2Plugin_logic_lq_regs_8_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_wordHit = ((Lsu2Plugin_logic_lq_regs_8_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_hit = ((((Lsu2Plugin_logic_lq_regs_8_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_wordHit) && Lsu2Plugin_logic_lq_regs_8_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[8]);
  assign when_Lsu2Plugin_l1104_8 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_8_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_pageHit = (Lsu2Plugin_logic_lq_regs_9_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_wordHit = ((Lsu2Plugin_logic_lq_regs_9_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_hit = ((((Lsu2Plugin_logic_lq_regs_9_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_wordHit) && Lsu2Plugin_logic_lq_regs_9_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[9]);
  assign when_Lsu2Plugin_l1104_9 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_9_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_pageHit = (Lsu2Plugin_logic_lq_regs_10_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_wordHit = ((Lsu2Plugin_logic_lq_regs_10_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_hit = ((((Lsu2Plugin_logic_lq_regs_10_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_wordHit) && Lsu2Plugin_logic_lq_regs_10_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[10]);
  assign when_Lsu2Plugin_l1104_10 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_10_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_pageHit = (Lsu2Plugin_logic_lq_regs_11_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_wordHit = ((Lsu2Plugin_logic_lq_regs_11_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_hit = ((((Lsu2Plugin_logic_lq_regs_11_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_wordHit) && Lsu2Plugin_logic_lq_regs_11_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[11]);
  assign when_Lsu2Plugin_l1104_11 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_11_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_pageHit = (Lsu2Plugin_logic_lq_regs_12_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_wordHit = ((Lsu2Plugin_logic_lq_regs_12_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_hit = ((((Lsu2Plugin_logic_lq_regs_12_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_wordHit) && Lsu2Plugin_logic_lq_regs_12_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[12]);
  assign when_Lsu2Plugin_l1104_12 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_12_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_pageHit = (Lsu2Plugin_logic_lq_regs_13_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_wordHit = ((Lsu2Plugin_logic_lq_regs_13_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_hit = ((((Lsu2Plugin_logic_lq_regs_13_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_wordHit) && Lsu2Plugin_logic_lq_regs_13_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[13]);
  assign when_Lsu2Plugin_l1104_13 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_13_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_pageHit = (Lsu2Plugin_logic_lq_regs_14_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_wordHit = ((Lsu2Plugin_logic_lq_regs_14_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_hit = ((((Lsu2Plugin_logic_lq_regs_14_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_wordHit) && Lsu2Plugin_logic_lq_regs_14_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[14]);
  assign when_Lsu2Plugin_l1104_14 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_14_hit);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_pageHit = (Lsu2Plugin_logic_lq_regs_15_address_pageOffset == Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 2]);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_wordHit = ((Lsu2Plugin_logic_lq_regs_15_address_mask & Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK) != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_hit = ((((Lsu2Plugin_logic_lq_regs_15_valid && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_pageHit) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_wordHit) && Lsu2Plugin_logic_lq_regs_15_sqChecked) && Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMask[15]);
  assign when_Lsu2Plugin_l1104_15 = ((! Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER) && Lsu2Plugin_logic_sharedPip_checkLqHits_entries_15_hit);
  assign Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER = Lsu2Plugin_logic_sharedPip_checkLqHits_youngerMaskEmpty;
  assign Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerHit = ((Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS != 16'h0000) && (! Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_NO_YOUNGER));
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_input = Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_priorityBits = Lsu2Plugin_logic_lq_ptr_priorityLast;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask = {Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_input,(Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_input[15 : 1] & Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_priorityBits)};
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 = Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[0];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_1 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[1];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[2];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[3];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[4];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_5 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[5];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[6];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_7 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[7];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[8];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[9];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[10];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_11 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[11];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[12];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_13 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[13];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_14 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[14];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_15 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[15];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_16 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[16];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_17 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[17];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_18 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[18];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_19 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[19];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_20 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[20];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_21 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[21];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_22 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[22];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_23 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[23];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_24 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[24];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_25 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[25];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_26 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[26];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_27 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[27];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_28 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[28];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_29 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[29];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_30 = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0[30];
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[0] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[1] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_1 && (! Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[2] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_2 && (! Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[3] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 && (! Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[4] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[5] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_5 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_4 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[6] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[7] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_7 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[8] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_8 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[9] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[10] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[11] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_11 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_10 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[12] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[13] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_13 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[14] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_14 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[15] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_15 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[16] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_16 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_15 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[17] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_17 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_16 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[18] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_18 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_17 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[19] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_19 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_18 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[20] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_20 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_19 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[21] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_21 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17)));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[22] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_22 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_21 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[23] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_23 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_22 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[24] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_24 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[25] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_25 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_24 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[26] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_26 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_25 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[27] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_27 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_26 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[28] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_28 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_27 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[29] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_29 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_28 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
    _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[30] = (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_30 && (! (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_29 || (Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26 || Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17))));
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_1 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_2,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_1,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_0}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_4 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_5,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_4,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_3}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_5 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_7 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_8,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_7,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_6}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_8 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_10 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_11,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_10,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_9}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_11 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2}}} != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_13 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_14,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_13,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_12}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_14 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2}}}} != 5'h00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_16 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_16,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_15} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_17 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_17,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_16,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_15}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_17 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_15_to_17,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_12_to_14,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_9_to_11,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_6_to_8,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_3_to_5,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_0_to_2}}}}} != 6'h00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_19 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_19,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_18} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_20,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_19,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_18}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_22 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_22,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_21} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_23,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_22,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_21}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_23 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_25 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_25,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_24} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_26 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_26,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_25,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_24}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_26 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_24_to_26,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_21_to_23,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_18_to_20}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_28 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_28,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_27} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_range_27_to_29 = ({Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_29,{Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_28,Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleMask_bools_27}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh = _zz_Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pLow = Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[30 : 15];
  assign Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pHigh = Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_doubleOh[14 : 0];
  assign Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh = (_zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh | Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS_roundRobinMasked_pLow);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[3];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_1 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[5];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_2 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[6];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[7];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_4 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[9];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_5 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[10];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_6 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[11];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_7 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[12];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_8 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[13];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_9 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[14];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_10 = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[15];
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_11 = (((((((Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[1] || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_1) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_4) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_6) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_8) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_10);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_12 = (((((((Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[2] || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_2) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_5) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_6) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_9) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_10);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_13 = (((((((Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[4] || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_1) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_2) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_3) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_7) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_8) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_9) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_10);
  assign _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_14 = (((((((Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerOh[8] || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_4) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_5) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_6) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_7) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_8) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_9) || _zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_10);
  assign Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel = {_zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_14,{_zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_13,{_zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_12,_zz_Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel_11}}};
  assign Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ROB = _zz_Lsu2Plugin_logic_lq_mem_robId_port2;
  assign Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_RESCHEDULE = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerHit;
  assign Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ID = Lsu2Plugin_logic_sharedPip_checkLqPrio_youngerSel;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride = 1'b1;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride = 1'b1;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_valid = Lsu2Plugin_setup_cacheLoad_rsp_valid;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data = Lsu2Plugin_setup_cacheLoad_rsp_payload_data;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data = LsuPlugin_peripheralBus_rsp_payload_data;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_fault = Lsu2Plugin_setup_cacheLoad_rsp_payload_fault;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_redo = Lsu2Plugin_setup_cacheLoad_rsp_payload_redo;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlot = Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlot;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlotAny = Lsu2Plugin_setup_cacheLoad_rsp_payload_refillSlotAny;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize = Lsu2Plugin_logic_sharedPip_stages_2_SIZE;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize = Lsu2Plugin_logic_special_loadSize;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize = Lsu2Plugin_logic_special_storeSize;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress = Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress = Lsu2Plugin_logic_special_loadAddress;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspAddress = Lsu2Plugin_logic_special_storeAddress;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned = Lsu2Plugin_logic_sharedPip_stages_2_UNSIGNED;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned = Lsu2Plugin_logic_special_loadUnsigned;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_0 = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data[7 : 0];
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_1 = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data[15 : 8];
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_2 = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data[23 : 16];
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3 = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data[31 : 24];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[7 : 0] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted;
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[15 : 8] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted_2;
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[23 : 16] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_2;
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[31 : 24] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspSplits_3;
    if(when_Lsu2Plugin_l1158) begin
      Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted = Lsu2Plugin_logic_sharedPip_checkSqArbi_bypass_data;
    end
  end

  assign when_Lsu2Plugin_l1158 = ((! Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride) && Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_HIT);
  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = (Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[7] && (! Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned));
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[31] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[30] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[29] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[28] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[27] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[26] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[25] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[24] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[23] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[22] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[21] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[20] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[19] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[18] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[17] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[16] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[15] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[14] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[13] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[12] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[11] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[10] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[9] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[8] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1[7 : 0] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[7 : 0];
  end

  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2 = (Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[15] && (! Lsu2Plugin_logic_sharedPip_cacheRsp_rspUnsigned));
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[31] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[30] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[29] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[28] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[27] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[26] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[25] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[24] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[23] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[22] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[21] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[20] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[19] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[18] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[17] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[16] = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_2;
    _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3[15 : 0] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[15 : 0];
  end

  assign _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_4[31 : 0] = Lsu2Plugin_logic_sharedPip_cacheRsp_rspShifted[31 : 0];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(Lsu2Plugin_logic_sharedPip_cacheRsp_rspSize)
      2'b00 : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_1;
      end
      2'b01 : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_3;
      end
      2'b10 : begin
        Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated = _zz_Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated_4;
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_isFireing = (Lsu2Plugin_logic_sharedPip_stages_2_valid && Lsu2Plugin_logic_sharedPip_stages_2_ready);
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_valid = ((Lsu2Plugin_logic_sharedPip_stages_2_isFireing && (! Lsu2Plugin_logic_sharedPip_stages_2_IS_IO)) && ((! Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION) || ((! Lsu2Plugin_logic_sharedPip_stages_2_MMU_REDO) && (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT))));
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_isLoad = Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_address = Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_TRANSLATED;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_readData = Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_robId = Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_lqId = Lsu2Plugin_logic_sharedPip_stages_2_LQ_ID;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_whitebox_size = Lsu2Plugin_logic_sharedPip_stages_2_SIZE;
  assign Lsu2Plugin_logic_sharedPip_cacheRsp_doIt = (((Lsu2Plugin_logic_sharedPip_stages_2_valid && Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD) && Lsu2Plugin_logic_sharedPip_stages_2_WRITE_RD) && ((! Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION) || ((Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_READ && (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT)) && (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_ACCESS_FAULT))));
  always @(*) begin
    Lsu2Plugin_setup_regfilePorts_0_write_valid = ((Lsu2Plugin_logic_sharedPip_cacheRsp_doIt && Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD) && 1'b1);
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_regfilePorts_0_write_valid = (Lsu2Plugin_logic_special_loadWriteRd && 1'b1);
    end
    if(Lsu2Plugin_logic_special_atomic_comp_rfWrite) begin
      Lsu2Plugin_setup_regfilePorts_0_write_valid = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_regfilePorts_0_write_address = Lsu2Plugin_logic_sharedPip_stages_2_PHYS_RD;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_regfilePorts_0_write_address = Lsu2Plugin_logic_special_loadPhysRd;
    end
    if(Lsu2Plugin_logic_special_atomic_comp_rfWrite) begin
      Lsu2Plugin_setup_regfilePorts_0_write_address = Lsu2Plugin_logic_sq_mem_physRd;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_regfilePorts_0_write_data = Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
        Lsu2Plugin_setup_regfilePorts_0_write_data = 32'h00000000;
        Lsu2Plugin_setup_regfilePorts_0_write_data[0] = (! Lsu2Plugin_logic_special_atomic_gotReservation);
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_regfilePorts_0_write_robId = Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_regfilePorts_0_write_robId = Lsu2Plugin_logic_special_robId;
    end
    if(Lsu2Plugin_logic_special_atomic_comp_rfWrite) begin
      Lsu2Plugin_setup_regfilePorts_0_write_robId = Lsu2Plugin_logic_special_robId;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_fpuWriteSize = Lsu2Plugin_logic_sharedPip_stages_2_SIZE;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_fpuWriteSize = Lsu2Plugin_logic_special_loadSize;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_WRITE_FAILURE = ((Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && Lsu2Plugin_logic_sharedPip_cacheRsp_specialOverride) && (! Lsu2Plugin_logic_sharedPip_stages_2_IS_IO));
  assign Lsu2Plugin_logic_sharedPip_stages_2_MISS_ALIGNED = ({((Lsu2Plugin_logic_sharedPip_stages_2_SIZE == 2'b10) && (Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION[1 : 0] != 2'b00)),((Lsu2Plugin_logic_sharedPip_stages_2_SIZE == 2'b01) && (Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION[0 : 0] != 1'b0))} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_stages_2_PAGE_FAULT = ((Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD ? (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_READ) : (! Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_WRITE)) || Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_cacheRsp_success = 1'b0;
    if(!Lsu2Plugin_logic_sharedPip_stages_2_MISS_ALIGNED) begin
      if(!when_Lsu2Plugin_l1203) begin
        if(!when_Lsu2Plugin_l1205) begin
          if(!when_Lsu2Plugin_l1207) begin
            if(!when_Lsu2Plugin_l1209) begin
              if(!when_Lsu2Plugin_l1211) begin
                if(!when_Lsu2Plugin_l1213) begin
                  Lsu2Plugin_logic_sharedPip_cacheRsp_success = 1'b1;
                end
              end
            end
          end
        end
      end
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_stages_2_MISS_ALIGNED) begin
      Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN;
    end else begin
      if(when_Lsu2Plugin_l1203) begin
        Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_MMU_REDO;
      end else begin
        if(when_Lsu2Plugin_l1205) begin
          Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_TRAP_MMU;
        end else begin
          if(when_Lsu2Plugin_l1207) begin
            Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD;
          end else begin
            if(when_Lsu2Plugin_l1209) begin
              Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_LOAD_MISS;
            end else begin
              if(when_Lsu2Plugin_l1211) begin
                Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_LOAD_FAILED;
              end else begin
                if(when_Lsu2Plugin_l1213) begin
                  Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS;
                end else begin
                  Lsu2Plugin_logic_sharedPip_stages_2_CTRL = Lsu2Plugin_CTRL_ENUM_SUCCESS;
                end
              end
            end
          end
        end
      end
    end
  end

  assign when_Lsu2Plugin_l1203 = (Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION && Lsu2Plugin_logic_sharedPip_stages_2_MMU_REDO);
  assign when_Lsu2Plugin_l1205 = (Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION && (Lsu2Plugin_logic_sharedPip_stages_2_MMU_ACCESS_FAULT || Lsu2Plugin_logic_sharedPip_stages_2_PAGE_FAULT));
  assign when_Lsu2Plugin_l1207 = (Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && ((Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_HIT && (! Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_BYPASS_SUCCESS)) || Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT));
  assign when_Lsu2Plugin_l1209 = (Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_redo);
  assign when_Lsu2Plugin_l1211 = (Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && Lsu2Plugin_logic_sharedPip_stages_2_LOAD_WRITE_FAILURE);
  assign when_Lsu2Plugin_l1213 = (Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD && Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_fault);
  assign Lsu2Plugin_logic_sharedPip_stages_2_TRAP_SPECULATION = (Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION && ((! Lsu2Plugin_logic_sharedPip_cacheRsp_success) || Lsu2Plugin_logic_sharedPip_stages_2_IS_IO));
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_valid = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_data = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_data;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_fault = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_fault;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_redo = Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_redo;
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny = (Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlotAny && (! (|DataCachePlugin_setup_refillCompletions)));
  assign Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlot = (Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_payload_refillSlot & (~ DataCachePlugin_setup_refillCompletions));
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_valid = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_data = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_data;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_fault = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_fault;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_redo = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_redo;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlotAny && (! (|DataCachePlugin_setup_refillCompletions)));
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlot = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlot & (~ DataCachePlugin_setup_refillCompletions));
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC = (Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD ? Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID : Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ID);
  assign Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC = _zz_Lsu2Plugin_logic_lq_mem_pc_port1;
  always @(*) begin
    Lsu2Plugin_setup_sharedCompletion_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(when_Lsu2Plugin_l1333) begin
              Lsu2Plugin_setup_sharedCompletion_valid = 1'b1;
            end
          end else begin
            if(when_Lsu2Plugin_l1374) begin
              Lsu2Plugin_setup_sharedCompletion_valid = 1'b1;
            end
          end
        end
      endcase
    end
  end

  assign Lsu2Plugin_setup_sharedCompletion_payload_id = Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(when_Lsu2Plugin_l1333) begin
              if(when_Lsu2Plugin_l1335) begin
                Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_valid = 1'b1;
              end
            end
          end
        end
      endcase
    end
  end

  assign Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_payload_robId = Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID;
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(when_Lsu2Plugin_l1333) begin
              if(when_Lsu2Plugin_l1335) begin
                Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid = 1'b1;
              end
            end
          end
        end
      endcase
    end
    if(Lsu2Plugin_logic_special_atomic_comp_wakeRf) begin
      Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_payload_physical = Lsu2Plugin_logic_sharedPip_stages_3_PHYS_RD;
    if(Lsu2Plugin_logic_special_atomic_comp_wakeRf) begin
      Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_payload_physical = Lsu2Plugin_logic_sq_mem_physRd;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_valid = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION) begin
        Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
      end
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
          Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
          Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
          Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_setup_sharedTrap_valid = 1'b1;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_payload_robId = Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_setup_sharedTrap_payload_robId = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ROB;
            end
          end
        end
      endcase
    end
  end

  assign Lsu2Plugin_setup_sharedTrap_payload_tval = Lsu2Plugin_logic_sharedPip_stages_3_ADDRESS_PRE_TRANSLATION;
  assign Lsu2Plugin_setup_sharedTrap_payload_skipCommit = 1'b1;
  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_payload_trap = 1'b1;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_setup_sharedTrap_payload_trap = 1'b0;
            end
          end
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_payload_cause = 4'bxxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION) begin
        Lsu2Plugin_setup_sharedTrap_payload_cause = 4'b1010;
      end
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
          Lsu2Plugin_setup_sharedTrap_payload_cause = 4'b0100;
          Lsu2Plugin_setup_sharedTrap_payload_cause[1] = (! Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD);
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
          Lsu2Plugin_setup_sharedTrap_payload_cause = 4'b1101;
          Lsu2Plugin_setup_sharedTrap_payload_cause[1] = (! Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD);
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
          Lsu2Plugin_setup_sharedTrap_payload_cause = 4'b0101;
          Lsu2Plugin_setup_sharedTrap_payload_cause[1] = (! Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_sharedTrap_payload_reason = 8'bxxxxxxxx;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      if(Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION) begin
        Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h03;
      end
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
          Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h01;
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
          Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h01;
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
          Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h01;
        end
        default : begin
          if(!Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE) begin
              Lsu2Plugin_setup_sharedTrap_payload_reason = 8'h20;
            end
          end
        end
      endcase
    end
  end

  assign Lsu2Plugin_setup_sharedTrap_payload_pcTarget = Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_PC;
  assign Lsu2Plugin_logic_sharedPip_ctrl_lqMask = (16'h0001 <<< Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID);
  assign Lsu2Plugin_logic_sharedPip_ctrl_sqMask = (16'h0001 <<< Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID);
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger = 1'b0;
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger = Lsu2Plugin_logic_translationWake;
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger = (! (|Lsu2Plugin_logic_sharedPip_ctrl_refillMask));
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
          Lsu2Plugin_logic_sharedPip_ctrl_redoTrigger = 1'b1;
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
        end
      endcase
    end
  end

  assign _zz_103 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[0];
  assign _zz_104 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[1];
  assign _zz_105 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[2];
  assign _zz_106 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[3];
  assign _zz_107 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[4];
  assign _zz_108 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[5];
  assign _zz_109 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[6];
  assign _zz_110 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[7];
  assign _zz_111 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[8];
  assign _zz_112 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[9];
  assign _zz_113 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[10];
  assign _zz_114 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[11];
  assign _zz_115 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[12];
  assign _zz_116 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[13];
  assign _zz_117 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[14];
  assign _zz_118 = Lsu2Plugin_logic_sharedPip_ctrl_lqMask[15];
  assign _zz_119 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[0];
  assign _zz_120 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[1];
  assign _zz_121 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[2];
  assign _zz_122 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[3];
  assign _zz_123 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[4];
  assign _zz_124 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[5];
  assign _zz_125 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[6];
  assign _zz_126 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[7];
  assign _zz_127 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[8];
  assign _zz_128 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[9];
  assign _zz_129 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[10];
  assign _zz_130 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[11];
  assign _zz_131 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[12];
  assign _zz_132 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[13];
  assign _zz_133 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[14];
  assign _zz_134 = Lsu2Plugin_logic_sharedPip_ctrl_sqMask[15];
  assign Lsu2Plugin_logic_sharedPip_ctrl_refillMask = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlotAny ? 2'b11 : Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlot);
  assign Lsu2Plugin_logic_sharedPip_ctrl_doCompletion = ((Lsu2Plugin_logic_sharedPip_stages_3_CTRL == Lsu2Plugin_CTRL_ENUM_SUCCESS) && (! Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION));
  assign Lsu2Plugin_logic_sharedPip_stages_3_isFireing = (Lsu2Plugin_logic_sharedPip_stages_3_valid && Lsu2Plugin_logic_sharedPip_stages_3_ready);
  assign when_Lsu2Plugin_l1313 = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT || Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_WAIT_FEED);
  assign _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT ? Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SQID : Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID);
  assign when_Lsu2Plugin_l1314 = (Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT ? Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_resulting : Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_resulting);
  assign when_Lsu2Plugin_l1333 = (! Lsu2Plugin_logic_sharedPip_stages_3_IS_IO);
  assign when_Lsu2Plugin_l1335 = (Lsu2Plugin_logic_sharedPip_stages_3_WRITE_RD && (! Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION));
  assign _zz_when_Lsu2Plugin_l1348 = _zz__zz_when_Lsu2Plugin_l1348;
  always @(*) begin
    _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'b000;
    if(when_Lsu2Plugin_l1348) begin
      _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'b001;
    end
    if(when_Lsu2Plugin_l1351) begin
      _zz_Lsu2Plugin_logic_lq_hazardPrediction_write_payload_data_score = 3'b111;
    end
  end

  assign when_Lsu2Plugin_l1348 = (_zz_when_Lsu2Plugin_l1348 && (&Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE));
  assign when_Lsu2Plugin_l1351 = ((! _zz_when_Lsu2Plugin_l1348) && (! (|Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE)));
  assign when_Lsu2Plugin_l1374 = (((! Lsu2Plugin_logic_sharedPip_stages_3_SC) && (! Lsu2Plugin_logic_sharedPip_stages_3_AMO)) && (! Lsu2Plugin_logic_sharedPip_stages_3_IS_IO));
  assign _zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next = ((Lsu2Plugin_logic_sharedPip_ctrl_doCompletion && (! Lsu2Plugin_logic_sharedPip_stages_3_IS_IO)) ? 6'h3f : 6'h14);
  assign Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next = ($signed(_zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_1) + $signed(_zz_Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next_2));
  assign Lsu2Plugin_logic_lq_hitPrediction_write_valid = (((Lsu2Plugin_logic_sharedPip_stages_3_isFireing && Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) && Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH) && (! Lsu2Plugin_logic_sharedPip_stages_3_SP_FP_ADDRESS));
  assign Lsu2Plugin_logic_lq_hitPrediction_write_payload_address = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH_PC[11 : 2];
  assign when_SInt_l131 = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[6];
  assign when_SInt_l132 = (! (&_zz_when_SInt_l132));
  always @(*) begin
    if(when_SInt_l131) begin
      if(when_SInt_l132) begin
        _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = 6'h20;
      end else begin
        _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[5 : 0];
      end
    end else begin
      if(when_SInt_l138) begin
        _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = 6'h1f;
      end else begin
        _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = Lsu2Plugin_logic_sharedPip_ctrl_hitPrediction_next[5 : 0];
      end
    end
  end

  assign when_SInt_l138 = (|_zz_when_SInt_l138);
  assign Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter = _zz_Lsu2Plugin_logic_lq_hitPrediction_write_payload_data_counter;
  assign Lsu2Plugin_logic_writeback_waitOn_ready = ((Lsu2Plugin_logic_writeback_waitOn_refillSlot == 2'b00) && (! Lsu2Plugin_logic_writeback_waitOn_refillSlotAny));
  always @(*) begin
    Lsu2Plugin_logic_writeback_waitOn_refillSlotSet = 2'b00;
    if(when_Lsu2Plugin_l1488) begin
      if(Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        Lsu2Plugin_logic_writeback_waitOn_refillSlotSet = Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlot;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_writeback_waitOn_refillSlotAnySet = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      if(Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        Lsu2Plugin_logic_writeback_waitOn_refillSlotAnySet = Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlotAny;
      end
    end
  end

  assign Lsu2Plugin_logic_writeback_feed_holdPrefetch = 1'b0;
  always @(*) begin
    Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready = toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready;
    if(when_Stream_l369_1) begin
      Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready = 1'b1;
    end
  end

  assign when_Stream_l369_1 = (! toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_valid);
  assign toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_valid = toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rValid;
  assign toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_payload = toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rData;
  assign _zz_toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready = (! Lsu2Plugin_logic_writeback_feed_holdPrefetch);
  assign toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready = (1'b1 && _zz_toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready);
  assign Lsu2Plugin_logic_writeback_feed_prediction_valid = (toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_valid && _zz_toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_ready);
  assign Lsu2Plugin_logic_writeback_feed_prediction_payload = toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_m2sPipe_payload;
  assign Lsu2Plugin_logic_writeback_feed_io = _zz_Lsu2Plugin_logic_sq_mem_io_port2[0];
  assign Lsu2Plugin_logic_writeback_feed_size = _zz_Lsu2Plugin_logic_sq_mem_size_port3;
  always @(*) begin
    Lsu2Plugin_logic_writeback_feed_data = _zz_Lsu2Plugin_logic_sq_mem_data_port2;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
        if(Lsu2Plugin_logic_special_storeAmo) begin
          Lsu2Plugin_logic_writeback_feed_data[31 : 0] = Lsu2Plugin_logic_special_atomic_result;
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_logic_writeback_feed_skip = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
        if(when_Lsu2Plugin_l1824) begin
          Lsu2Plugin_logic_writeback_feed_skip = 1'b1;
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_writeback_feed_doit = (((Lsu2Plugin_logic_sq_ptr_writeBack != Lsu2Plugin_logic_sq_ptr_commit) && Lsu2Plugin_logic_writeback_waitOn_ready) && (! Lsu2Plugin_logic_writeback_feed_prediction_valid));
  always @(*) begin
    Lsu2Plugin_logic_writeback_feed_fire = (Lsu2Plugin_logic_writeback_feed_doit && Lsu2Plugin_setup_cacheStore_cmd_ready);
    if(when_Lsu2Plugin_l1509) begin
      Lsu2Plugin_logic_writeback_feed_fire = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_valid = Lsu2Plugin_logic_writeback_feed_doit;
    if(Lsu2Plugin_logic_writeback_feed_prediction_valid) begin
      Lsu2Plugin_setup_cacheStore_cmd_valid = 1'b1;
    end
    if(when_Lsu2Plugin_l1509) begin
      Lsu2Plugin_setup_cacheStore_cmd_valid = 1'b0;
    end
    if(when_Lsu2Plugin_l1553) begin
      Lsu2Plugin_setup_cacheStore_cmd_valid = (! Lsu2Plugin_logic_flush_cmdPtr[6]);
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_address = _zz_Lsu2Plugin_logic_sq_mem_addressPost_port3;
    if(Lsu2Plugin_logic_writeback_feed_prediction_valid) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_address = Lsu2Plugin_logic_writeback_feed_prediction_payload;
    end
    if(when_Lsu2Plugin_l1553) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_address[11 : 6] = Lsu2Plugin_logic_flush_cmdPtr[5:0];
    end
  end

  always @(*) begin
    _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask = 4'bxxxx;
    case(Lsu2Plugin_logic_writeback_feed_size)
      2'b00 : begin
        _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask = 4'b0001;
      end
      2'b01 : begin
        _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask = 4'b0011;
      end
      2'b10 : begin
        _zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask = 4'b1111;
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_cacheStore_cmd_payload_mask = (_zz_Lsu2Plugin_setup_cacheStore_cmd_payload_mask <<< Lsu2Plugin_setup_cacheStore_cmd_payload_address[1 : 0]);
  assign Lsu2Plugin_setup_cacheStore_cmd_payload_generation = Lsu2Plugin_logic_writeback_generation;
  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(Lsu2Plugin_logic_writeback_feed_size)
      2'b00 : begin
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[7 : 0] = Lsu2Plugin_logic_writeback_feed_data[7 : 0];
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[15 : 8] = Lsu2Plugin_logic_writeback_feed_data[7 : 0];
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[23 : 16] = Lsu2Plugin_logic_writeback_feed_data[7 : 0];
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[31 : 24] = Lsu2Plugin_logic_writeback_feed_data[7 : 0];
      end
      2'b01 : begin
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[15 : 0] = Lsu2Plugin_logic_writeback_feed_data[15 : 0];
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[31 : 16] = Lsu2Plugin_logic_writeback_feed_data[15 : 0];
      end
      2'b10 : begin
        Lsu2Plugin_setup_cacheStore_cmd_payload_data[31 : 0] = Lsu2Plugin_logic_writeback_feed_data[31 : 0];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_io = Lsu2Plugin_logic_writeback_feed_io;
    if(Lsu2Plugin_logic_writeback_feed_prediction_valid) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_io = 1'b0;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_prefetch = 1'b0;
    if(Lsu2Plugin_logic_writeback_feed_prediction_valid) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_prefetch = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_valid = Lsu2Plugin_setup_cacheStore_rsp_valid;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_fault = Lsu2Plugin_setup_cacheStore_rsp_payload_fault;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_redo = Lsu2Plugin_setup_cacheStore_rsp_payload_redo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlot = Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlot;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlotAny = Lsu2Plugin_setup_cacheStore_rsp_payload_refillSlotAny;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_generationKo = Lsu2Plugin_setup_cacheStore_rsp_payload_generationKo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_flush = Lsu2Plugin_setup_cacheStore_rsp_payload_flush;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_prefetch = Lsu2Plugin_setup_cacheStore_rsp_payload_prefetch;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_address = Lsu2Plugin_setup_cacheStore_rsp_payload_address;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_io = Lsu2Plugin_setup_cacheStore_rsp_payload_io;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_valid = Lsu2Plugin_logic_writeback_rsp_delayed_0_valid;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_fault = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_fault;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_redo = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_redo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_generationKo = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_generationKo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_flush = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_flush;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_prefetch = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_prefetch;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_address = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_address;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_io = Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_io;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_valid = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_valid;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_fault = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_fault;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_redo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlot = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlot;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlotAny = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlotAny;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_generationKo = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_generationKo;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_flush = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_flush;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_prefetch = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_prefetch;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_address = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_address;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_io = Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_io;
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlot = (Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlot & (~ DataCachePlugin_setup_refillCompletions));
  assign Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlotAny = (Lsu2Plugin_logic_writeback_rsp_delayed_0_payload_refillSlotAny && (DataCachePlugin_setup_refillCompletions == 2'b00));
  always @(*) begin
    Lsu2Plugin_logic_sq_ptr_onFree_valid = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      if(!Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        Lsu2Plugin_logic_sq_ptr_onFree_valid = 1'b1;
      end
    end
    if(when_Lsu2Plugin_l1509) begin
      Lsu2Plugin_logic_sq_ptr_onFree_valid = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_sq_ptr_onFree_payload = Lsu2Plugin_logic_sq_ptr_freeReal;
  always @(*) begin
    Lsu2Plugin_logic_writeback_rsp_whitebox_valid = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      if(!Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        if(when_Lsu2Plugin_l1498) begin
          Lsu2Plugin_logic_writeback_rsp_whitebox_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_prefetch_predictor_io_learn_valid = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      Lsu2Plugin_logic_prefetch_predictor_io_learn_valid = 1'b1;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_prefetch_predictor_io_learn_payload_allocate = 1'b0;
    if(when_Lsu2Plugin_l1488) begin
      if(Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
        Lsu2Plugin_logic_prefetch_predictor_io_learn_payload_allocate = 1'b1;
      end
    end
  end

  assign when_Lsu2Plugin_l1488 = (((Lsu2Plugin_logic_writeback_rsp_delayed_1_valid && (! Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_generationKo)) && (! Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_flush)) && (! Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_prefetch));
  assign when_Lsu2Plugin_l1498 = (! Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_io);
  assign Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_valid = (Lsu2Plugin_logic_writeback_rsp_delayed_1_valid && Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_prefetch);
  assign Lsu2Plugin_logic_prefetch_predictor_io_prediction_rsp_payload = (|Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_refillSlot);
  assign when_Lsu2Plugin_l1509 = (Lsu2Plugin_logic_writeback_feed_doit && Lsu2Plugin_logic_writeback_feed_skip);
  always @(*) begin
    Lsu2Plugin_logic_sq_tracker_add = 1'b0;
    if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
      Lsu2Plugin_logic_sq_tracker_add = 1'b1;
    end
  end

  assign when_Lsu2Plugin_l1521 = (Lsu2Plugin_logic_sq_ptr_priority == 15'h0000);
  assign when_Lsu2Plugin_l1524 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b0000);
  assign when_Lsu2Plugin_l1524_1 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b0001);
  assign when_Lsu2Plugin_l1524_2 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b0010);
  assign when_Lsu2Plugin_l1524_3 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b0011);
  assign when_Lsu2Plugin_l1524_4 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b0100);
  assign when_Lsu2Plugin_l1524_5 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b0101);
  assign when_Lsu2Plugin_l1524_6 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b0110);
  assign when_Lsu2Plugin_l1524_7 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b0111);
  assign when_Lsu2Plugin_l1524_8 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b1000);
  assign when_Lsu2Plugin_l1524_9 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b1001);
  assign when_Lsu2Plugin_l1524_10 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b1010);
  assign when_Lsu2Plugin_l1524_11 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b1011);
  assign when_Lsu2Plugin_l1524_12 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b1100);
  assign when_Lsu2Plugin_l1524_13 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b1101);
  assign when_Lsu2Plugin_l1524_14 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b1110);
  assign when_Lsu2Plugin_l1524_15 = (Lsu2Plugin_logic_sq_ptr_freeReal == 4'b1111);
  assign FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548 = _zz_FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548;
  always @(*) begin
    Lsu2Plugin_setup_cacheStore_cmd_payload_flush = 1'b0;
    if(when_Lsu2Plugin_l1553) begin
      Lsu2Plugin_setup_cacheStore_cmd_payload_flush = 1'b1;
    end
  end

  assign Lsu2Plugin_setup_cacheStore_cmd_payload_flushFree = Lsu2Plugin_logic_flush_withFree;
  assign when_Lsu2Plugin_l1553 = (Lsu2Plugin_logic_flush_busy && Lsu2Plugin_logic_flush_doit);
  assign Lsu2Plugin_setup_cacheStore_cmd_fire = (Lsu2Plugin_setup_cacheStore_cmd_valid && Lsu2Plugin_setup_cacheStore_cmd_ready);
  assign when_Lsu2Plugin_l1561 = (Lsu2Plugin_setup_cacheStore_rsp_valid && (! Lsu2Plugin_setup_cacheStore_rsp_payload_generationKo));
  assign when_Lsu2Plugin_l1569 = (Lsu2Plugin_logic_flush_rspPtr[6] && (! DataCachePlugin_setup_writebackBusy));
  assign Lsu2Plugin_logic_special_lqOnTop = (_zz_Lsu2Plugin_logic_lq_mem_robId_port3 == CommitPlugin_logic_commit_head);
  assign Lsu2Plugin_logic_special_sqOnTop = (_zz_Lsu2Plugin_logic_sq_mem_robId_port2 == CommitPlugin_logic_commit_head);
  assign Lsu2Plugin_logic_special_storeWriteBackUsable = (Lsu2Plugin_logic_sq_ptr_writeBack == Lsu2Plugin_logic_sq_ptr_commit);
  assign Lsu2Plugin_logic_special_storeSpecial = Lsu2Plugin_logic_sq_mem_doSpecial_io_read_0_rsp[0];
  assign Lsu2Plugin_logic_special_loadSpecial = Lsu2Plugin_logic_lq_mem_doSpecial_io_read_0_rsp[0];
  assign Lsu2Plugin_logic_special_storeHit = (((Lsu2Plugin_logic_special_sqOnTop && Lsu2Plugin_logic_special_storeWriteBackUsable) && (Lsu2Plugin_logic_sq_ptr_commit != Lsu2Plugin_logic_sq_ptr_alloc)) && Lsu2Plugin_logic_special_storeSpecial);
  assign Lsu2Plugin_logic_special_loadHit = ((Lsu2Plugin_logic_special_lqOnTop && (Lsu2Plugin_logic_lq_ptr_free != Lsu2Plugin_logic_lq_ptr_alloc)) && Lsu2Plugin_logic_special_loadSpecial);
  assign Lsu2Plugin_logic_special_hit = (Lsu2Plugin_logic_special_storeHit || Lsu2Plugin_logic_special_loadHit);
  always @(*) begin
    Lsu2Plugin_logic_special_fire = LsuPlugin_peripheralBus_rsp_valid_regNext;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
        if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
          Lsu2Plugin_logic_special_fire = 1'b1;
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  assign LsuPlugin_peripheralBus_cmd_fire = (LsuPlugin_peripheralBus_cmd_valid && LsuPlugin_peripheralBus_cmd_ready);
  assign Lsu2Plugin_logic_special_address = (Lsu2Plugin_logic_special_isStore ? Lsu2Plugin_logic_special_storeAddress : Lsu2Plugin_logic_special_loadAddress);
  assign Lsu2Plugin_logic_special_addressVirt = (Lsu2Plugin_logic_special_isStore ? Lsu2Plugin_logic_special_storeAddressVirt : Lsu2Plugin_logic_special_loadAddressVirt);
  assign Lsu2Plugin_logic_special_isIo = (! (Lsu2Plugin_logic_special_isStore && (Lsu2Plugin_logic_special_storeAmo || Lsu2Plugin_logic_special_storeSc)));
  assign Lsu2Plugin_logic_special_isAtomic = (! Lsu2Plugin_logic_special_isIo);
  always @(*) begin
    Lsu2Plugin_logic_special_wakeRob_valid = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      if(Lsu2Plugin_logic_special_loadWriteRd) begin
        Lsu2Plugin_logic_special_wakeRob_valid = 1'b1;
      end
    end
    if(Lsu2Plugin_logic_special_atomic_comp_wakeRf) begin
      Lsu2Plugin_logic_special_wakeRob_valid = 1'b1;
    end
  end

  assign Lsu2Plugin_logic_special_wakeRob_payload_robId = Lsu2Plugin_logic_special_robId;
  always @(*) begin
    Lsu2Plugin_logic_special_wakeRf_valid = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      if(Lsu2Plugin_logic_special_loadWriteRd) begin
        Lsu2Plugin_logic_special_wakeRf_valid = 1'b1;
      end
    end
  end

  assign Lsu2Plugin_logic_special_wakeRf_payload_physical = Lsu2Plugin_logic_special_loadPhysRd;
  assign LsuPlugin_peripheralBus_cmd_valid = ((Lsu2Plugin_logic_special_enabled && (! Lsu2Plugin_logic_special_cmdSent)) && Lsu2Plugin_logic_special_isIo);
  assign LsuPlugin_peripheralBus_cmd_payload_write = Lsu2Plugin_logic_special_isStore;
  assign LsuPlugin_peripheralBus_cmd_payload_address = Lsu2Plugin_logic_special_address;
  assign LsuPlugin_peripheralBus_cmd_payload_size = (Lsu2Plugin_logic_special_isStore ? Lsu2Plugin_logic_special_storeSize : Lsu2Plugin_logic_special_loadSize);
  assign LsuPlugin_peripheralBus_cmd_payload_data = Lsu2Plugin_logic_special_storeData;
  assign LsuPlugin_peripheralBus_cmd_payload_mask = Lsu2Plugin_logic_special_storeMask;
  always @(*) begin
    Lsu2Plugin_setup_specialTrap_valid = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_specialTrap_valid = LsuPlugin_peripheralBus_rsp_payload_error;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
        Lsu2Plugin_setup_specialTrap_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_specialTrap_payload_robId = Lsu2Plugin_logic_special_robId;
  assign Lsu2Plugin_setup_specialTrap_payload_cause = {1'd0, _zz_Lsu2Plugin_setup_specialTrap_payload_cause};
  assign Lsu2Plugin_setup_specialTrap_payload_tval = Lsu2Plugin_logic_special_addressVirt;
  assign Lsu2Plugin_setup_specialTrap_payload_skipCommit = 1'b1;
  assign Lsu2Plugin_setup_specialTrap_payload_reason = 8'h01;
  always @(*) begin
    Lsu2Plugin_setup_specialCompletion_valid = 1'b0;
    if(LsuPlugin_peripheralBus_rsp_valid) begin
      Lsu2Plugin_setup_specialCompletion_valid = 1'b1;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
        Lsu2Plugin_setup_specialCompletion_valid = 1'b1;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_specialCompletion_payload_id = Lsu2Plugin_logic_special_robId;
  assign Lsu2Plugin_logic_special_atomic_wantExit = 1'b0;
  always @(*) begin
    Lsu2Plugin_logic_special_atomic_wantStart = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
        Lsu2Plugin_logic_special_atomic_wantStart = 1'b1;
      end
    endcase
  end

  assign Lsu2Plugin_logic_special_atomic_wantKill = 1'b0;
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub = Lsu2Plugin_logic_special_atomic_readed[31 : 0];
  assign _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 = Lsu2Plugin_logic_special_storeData[31 : 0];
  assign Lsu2Plugin_logic_special_atomic_alu_compare = Lsu2Plugin_logic_sq_mem_op[2];
  assign Lsu2Plugin_logic_special_atomic_alu_unsigned = Lsu2Plugin_logic_sq_mem_op[1];
  assign Lsu2Plugin_logic_special_atomic_alu_addSub = _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_2;
  assign Lsu2Plugin_logic_special_atomic_alu_less = ((_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1[31] == _zz_Lsu2Plugin_logic_special_atomic_alu_addSub[31]) ? Lsu2Plugin_logic_special_atomic_alu_addSub[31] : (Lsu2Plugin_logic_special_atomic_alu_unsigned ? _zz_Lsu2Plugin_logic_special_atomic_alu_addSub[31] : _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1[31]));
  assign Lsu2Plugin_logic_special_atomic_alu_selectRf = (Lsu2Plugin_logic_sq_mem_swap ? 1'b1 : (Lsu2Plugin_logic_sq_mem_op[0] ^ Lsu2Plugin_logic_special_atomic_alu_less));
  assign switch_Misc_l232_2 = (Lsu2Plugin_logic_sq_mem_op | {Lsu2Plugin_logic_sq_mem_swap,2'b00});
  always @(*) begin
    case(switch_Misc_l232_2)
      3'b000 : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = Lsu2Plugin_logic_special_atomic_alu_addSub;
      end
      3'b001 : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = (_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 ^ _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
      end
      3'b010 : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = (_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 | _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
      end
      3'b011 : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = (_zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 & _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
      end
      default : begin
        Lsu2Plugin_logic_special_atomic_alu_raw = (Lsu2Plugin_logic_special_atomic_alu_selectRf ? _zz_Lsu2Plugin_logic_special_atomic_alu_addSub_1 : _zz_Lsu2Plugin_logic_special_atomic_alu_addSub);
      end
    endcase
  end

  assign Lsu2Plugin_logic_special_atomic_alu_result = Lsu2Plugin_logic_special_atomic_alu_raw;
  assign when_Lsu2Plugin_l1683 = (Lsu2Plugin_logic_special_enabled && Lsu2Plugin_logic_special_isAtomic);
  always @(*) begin
    DataCachePlugin_setup_lockPort_valid = 1'b0;
    if(when_Lsu2Plugin_l1698) begin
      DataCachePlugin_setup_lockPort_valid = 1'b1;
    end
  end

  always @(*) begin
    DataCachePlugin_setup_lockPort_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_Lsu2Plugin_l1698) begin
      DataCachePlugin_setup_lockPort_address = Lsu2Plugin_logic_special_storeAddress;
    end
  end

  assign Lsu2Plugin_setup_cacheLoad_cmd_payload_unlocked = 1'b1;
  assign when_Lsu2Plugin_l1698 = (! ((Lsu2Plugin_logic_special_atomic_stateReg & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) != 9'b000000000));
  always @(*) begin
    Lsu2Plugin_logic_special_atomic_loadWhitebox_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
        if(Lsu2Plugin_setup_cacheLoad_rsp_valid) begin
          if(!Lsu2Plugin_setup_cacheLoad_rsp_payload_redo) begin
            if(!Lsu2Plugin_setup_cacheLoad_rsp_payload_fault) begin
              Lsu2Plugin_logic_special_atomic_loadWhitebox_valid = 1'b1;
            end
          end
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_special_atomic_loadWhitebox_readData = Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated[31 : 0];
  always @(*) begin
    Lsu2Plugin_logic_special_atomic_storeWhitebox_valid = 1'b0;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
        Lsu2Plugin_logic_special_atomic_storeWhitebox_valid = 1'b1;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_logic_special_atomic_storeWhitebox_isSc = Lsu2Plugin_logic_special_storeSc;
  assign Lsu2Plugin_logic_special_atomic_storeWhitebox_scPassed = Lsu2Plugin_logic_special_atomic_gotReservation;
  assign FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l1834 = ((Lsu2Plugin_logic_special_atomic_stateReg & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) != 9'b000000000);
  always @(*) begin
    Lsu2Plugin_logic_lqFlush = 1'b0;
    if(CommitPlugin_logic_commit_reschedulePort_valid) begin
      Lsu2Plugin_logic_lqFlush = 1'b1;
    end
  end

  assign when_Lsu2Plugin_l1909 = (! Lsu2Plugin_logic_sq_regs_0_commitedNext);
  assign when_Lsu2Plugin_l1909_1 = (! Lsu2Plugin_logic_sq_regs_1_commitedNext);
  assign when_Lsu2Plugin_l1909_2 = (! Lsu2Plugin_logic_sq_regs_2_commitedNext);
  assign when_Lsu2Plugin_l1909_3 = (! Lsu2Plugin_logic_sq_regs_3_commitedNext);
  assign when_Lsu2Plugin_l1909_4 = (! Lsu2Plugin_logic_sq_regs_4_commitedNext);
  assign when_Lsu2Plugin_l1909_5 = (! Lsu2Plugin_logic_sq_regs_5_commitedNext);
  assign when_Lsu2Plugin_l1909_6 = (! Lsu2Plugin_logic_sq_regs_6_commitedNext);
  assign when_Lsu2Plugin_l1909_7 = (! Lsu2Plugin_logic_sq_regs_7_commitedNext);
  assign when_Lsu2Plugin_l1909_8 = (! Lsu2Plugin_logic_sq_regs_8_commitedNext);
  assign when_Lsu2Plugin_l1909_9 = (! Lsu2Plugin_logic_sq_regs_9_commitedNext);
  assign when_Lsu2Plugin_l1909_10 = (! Lsu2Plugin_logic_sq_regs_10_commitedNext);
  assign when_Lsu2Plugin_l1909_11 = (! Lsu2Plugin_logic_sq_regs_11_commitedNext);
  assign when_Lsu2Plugin_l1909_12 = (! Lsu2Plugin_logic_sq_regs_12_commitedNext);
  assign when_Lsu2Plugin_l1909_13 = (! Lsu2Plugin_logic_sq_regs_13_commitedNext);
  assign when_Lsu2Plugin_l1909_14 = (! Lsu2Plugin_logic_sq_regs_14_commitedNext);
  assign when_Lsu2Plugin_l1909_15 = (! Lsu2Plugin_logic_sq_regs_15_commitedNext);
  assign sqAlloc_0_valid = ((FrontendPlugin_dispatch_isFireing && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && FrontendPlugin_dispatch_SQ_ALLOC_0);
  assign sqAlloc_0_id = FrontendPlugin_dispatch_SQ_ID_0;
  assign sqAlloc_1_valid = ((FrontendPlugin_dispatch_isFireing && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1) && FrontendPlugin_dispatch_SQ_ALLOC_1);
  assign sqAlloc_1_id = FrontendPlugin_dispatch_SQ_ID_1;
  assign sqFree_valid = Lsu2Plugin_logic_sq_ptr_onFree_valid;
  assign sqFree_payload = Lsu2Plugin_logic_sq_ptr_onFree_payload;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken = BranchContextPlugin_logic_mem_earlyBranch_io_read_0_rsp;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken = _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken[0];
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc = _zz_ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken[32 : 1];
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BAD_EARLY_TARGET = (ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc != ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE);
  assign ALU0_BranchPlugin_setup_intFormatPort_payload = _zz_ALU0_BranchPlugin_setup_intFormatPort_payload;
  assign ALU0_BranchPlugin_logic_branch_badEarlyTaken = (ALU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_taken != ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND);
  assign ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSPREDICTED = (ALU0_BranchPlugin_logic_branch_badEarlyTaken || (ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND && ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BAD_EARLY_TARGET));
  assign ALU0_BranchPlugin_setup_reschedule_payload_robId = ALU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
  assign ALU0_BranchPlugin_setup_reschedule_payload_pcTarget = ALU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET;
  assign ALU0_BranchPlugin_setup_reschedule_payload_reason = {3'd0, _zz_ALU0_BranchPlugin_setup_reschedule_payload_reason};
  assign ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED = ((ALU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET[1 : 0] != 2'b00) && ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND);
  assign ALU0_ExecutionUnitBase_pipeline_execute_1_isFireing = (ALU0_ExecutionUnitBase_pipeline_execute_1_valid && ALU0_ExecutionUnitBase_pipeline_execute_1_ready);
  assign ALU0_BranchPlugin_setup_reschedule_valid = ((ALU0_ExecutionUnitBase_pipeline_execute_1_isFireing && ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL) && (ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSPREDICTED || ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED));
  assign ALU0_BranchPlugin_setup_reschedule_payload_trap = ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED;
  assign ALU0_BranchPlugin_setup_reschedule_payload_skipCommit = ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED;
  assign ALU0_BranchPlugin_setup_reschedule_payload_cause = 4'b0000;
  assign ALU0_BranchPlugin_setup_reschedule_payload_tval = ALU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET;
  assign ALU0_BranchPlugin_logic_branch_finalBranch_valid = (ALU0_ExecutionUnitBase_pipeline_execute_1_valid && ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL);
  assign ALU0_BranchPlugin_logic_branch_finalBranch_payload_address = ALU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_ID;
  assign ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice = (ALU0_ExecutionUnitBase_pipeline_execute_1_PC + _zz_ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice);
  assign ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcTarget = ALU0_ExecutionUnitBase_pipeline_execute_1_PC_TRUE;
  assign ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_taken = ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND;
  assign _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken = BranchContextPlugin_logic_mem_earlyBranch_io_read_1_rsp;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken = _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken[0];
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc = _zz_ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken[32 : 1];
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BAD_EARLY_TARGET = (ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc != ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TRUE);
  assign ALU1_BranchPlugin_setup_intFormatPort_payload = _zz_ALU1_BranchPlugin_setup_intFormatPort_payload;
  assign ALU1_BranchPlugin_logic_branch_badEarlyTaken = (ALU1_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_taken != ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND);
  assign ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSPREDICTED = (ALU1_BranchPlugin_logic_branch_badEarlyTaken || (ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND && ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BAD_EARLY_TARGET));
  assign ALU1_BranchPlugin_setup_reschedule_payload_robId = ALU1_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
  assign ALU1_BranchPlugin_setup_reschedule_payload_pcTarget = ALU1_ExecutionUnitBase_pipeline_execute_1_PC_TARGET;
  assign ALU1_BranchPlugin_setup_reschedule_payload_reason = {3'd0, _zz_ALU1_BranchPlugin_setup_reschedule_payload_reason};
  assign ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED = ((ALU1_ExecutionUnitBase_pipeline_execute_1_PC_TARGET[1 : 0] != 2'b00) && ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND);
  assign ALU1_ExecutionUnitBase_pipeline_execute_1_isFireing = (ALU1_ExecutionUnitBase_pipeline_execute_1_valid && ALU1_ExecutionUnitBase_pipeline_execute_1_ready);
  assign ALU1_BranchPlugin_setup_reschedule_valid = ((ALU1_ExecutionUnitBase_pipeline_execute_1_isFireing && ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL) && (ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSPREDICTED || ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED));
  assign ALU1_BranchPlugin_setup_reschedule_payload_trap = ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED;
  assign ALU1_BranchPlugin_setup_reschedule_payload_skipCommit = ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_MISSALIGNED;
  assign ALU1_BranchPlugin_setup_reschedule_payload_cause = 4'b0000;
  assign ALU1_BranchPlugin_setup_reschedule_payload_tval = ALU1_ExecutionUnitBase_pipeline_execute_1_PC_TARGET;
  assign ALU1_BranchPlugin_logic_branch_finalBranch_valid = (ALU1_ExecutionUnitBase_pipeline_execute_1_valid && ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL);
  assign ALU1_BranchPlugin_logic_branch_finalBranch_payload_address = ALU1_ExecutionUnitBase_pipeline_execute_1_BRANCH_ID;
  assign ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice = (ALU1_ExecutionUnitBase_pipeline_execute_1_PC + _zz_ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice);
  assign ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcTarget = ALU1_ExecutionUnitBase_pipeline_execute_1_PC_TRUE;
  assign ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_taken = ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND;
  assign MmuPlugin_logic_satpModeWrite = EU0_CsrAccessPlugin_setup_onWriteBits[31 : 31];
  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_refillOngoing = 1'b0;
    if(MmuPlugin_logic_refill_busy) begin
      if(_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask) begin
        FetchCachePlugin_setup_translationStorage_logic_refillOngoing = 1'b1;
      end
    end
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask = 4'b0000;
    if(when_MmuPlugin_l492) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask = 4'b1111;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask = ((_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask != 1'b0) ? _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask_1 : 4'b0000);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address = 5'bxxxxx;
    if(when_MmuPlugin_l492) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter[4:0];
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[16 : 12];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(when_MmuPlugin_l492) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_0) || (! MmuPlugin_logic_refill_load_flags_A));
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_accessFault = ((! FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_pageFault) && 1'b0);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress = 15'bxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 17];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value == 2'b11);
  assign FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflow = (FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc && FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext = (FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value + _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext);
    if(FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_willClear) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext = 2'b00;
    end
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask = 2'b00;
    if(when_MmuPlugin_l492) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask = 2'b11;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask = ((_zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask != 1'b0) ? _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_write_mask : 2'b00);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address = 5'bxxxxx;
    if(when_MmuPlugin_l492) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter[4:0];
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[26 : 22];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(when_MmuPlugin_l492) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_1) || (! MmuPlugin_logic_refill_load_flags_A));
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_accessFault = ((! FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_pageFault) && 1'b0);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress = 5'bxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 27];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress = 10'bxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd22);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc = (FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value == 1'b1);
  assign FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflow = (FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc && FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement);
  always @(*) begin
    FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_valueNext = (FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value + FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willIncrement);
    if(FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_willClear) begin
      FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_valueNext = 1'b0;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_refillOngoing = 1'b0;
    if(MmuPlugin_logic_refill_busy) begin
      if(_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask) begin
        Lsu2Plugin_setup_translationStorage_logic_refillOngoing = 1'b1;
      end
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask = 4'b0000;
    if(when_MmuPlugin_l492) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask = 4'b1111;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask = ((_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask != 1'b0) ? _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask_1 : 4'b0000);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address = 5'bxxxxx;
    if(when_MmuPlugin_l492) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter[4:0];
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[16 : 12];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(when_MmuPlugin_l492) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_valid = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_0) || (! MmuPlugin_logic_refill_load_flags_A));
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_accessFault = ((! Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_pageFault) && 1'b0);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress = 15'bxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 17];
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value == 2'b11);
  assign Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflow = (Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willOverflowIfInc && Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext = (Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value + _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext);
    if(Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_willClear) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext = 2'b00;
    end
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask = 2'b00;
    if(when_MmuPlugin_l492) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask = 2'b11;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask = ((_zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask != 1'b0) ? _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_write_mask : 2'b00);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address = 5'bxxxxx;
    if(when_MmuPlugin_l492) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter[4:0];
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[26 : 22];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(when_MmuPlugin_l492) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_valid = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_1) || (! MmuPlugin_logic_refill_load_flags_A));
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_accessFault = ((! Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_pageFault) && 1'b0);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress = 5'bxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 27];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress = 10'bxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd22);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l469) begin
              Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc = (Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value == 1'b1);
  assign Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflow = (Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willOverflowIfInc && Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement);
  always @(*) begin
    Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_valueNext = (Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value + Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willIncrement);
    if(Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_willClear) begin
      Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_valueNext = 1'b0;
    end
  end

  assign Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL = Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL_overloaded = ((Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL && (! Lsu2Plugin_setup_translationStorage_logic_refillOngoing)) && Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg);
  assign when_MmuPlugin_l260 = (Lsu2Plugin_logic_sharedPip_stages_0_isRemoved || (! (Lsu2Plugin_logic_sharedPip_stages_0_valid && (! Lsu2Plugin_logic_sharedPip_stages_0_ready))));
  assign Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded = ((Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL && (! Lsu2Plugin_setup_translationStorage_logic_refillOngoing)) && Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg);
  assign when_MmuPlugin_l260_1 = (Lsu2Plugin_logic_sharedPip_stages_1_isRemoved || (! (Lsu2Plugin_logic_sharedPip_stages_1_valid && (! Lsu2Plugin_logic_sharedPip_stages_1_ready))));
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_read_0_readAddress = Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[16 : 12];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid = _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_0_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[17 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[37 : 18];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[38];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[39];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[40];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid[41];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID[0] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 17]);
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID[1] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 17]);
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID[2] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 17]);
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID[3] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 17]);
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS[0] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID[0] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_valid);
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS[1] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID[1] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_valid);
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS[2] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID[2] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_valid);
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS[3] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID[3] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_valid);
  end

  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid = _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_1_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[17 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[37 : 18];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[38];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[39];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[40];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid[41];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid = _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_2_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[17 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[37 : 18];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[38];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[39];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[40];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid[41];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid = _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_ways_3_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[17 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[37 : 18];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[38];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[39];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[40];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid[41];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_read_1_readAddress = Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[26 : 22];
  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid = _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_0_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[7 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[17 : 8];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[18];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[19];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[20];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid[21];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_HITS_PRE_VALID[0] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 27]);
    Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_HITS_PRE_VALID[1] = (Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_virtualAddress == Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION[31 : 27]);
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS[0] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS_PRE_VALID[0] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_valid);
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS[1] = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS_PRE_VALID[1] && Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_valid);
  end

  assign _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid = _zz_Lsu2Plugin_setup_translationStorage_logic_sl_1_ways_1_port1;
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[0];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_pageFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[1];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_accessFault = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[2];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_virtualAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[7 : 3];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_physicalAddress = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[17 : 8];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowRead = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[18];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowWrite = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[19];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowExecute = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[20];
  assign Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowUser = _zz_Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid[21];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS,Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS};
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hit = (|Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits);
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits;
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[1];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[2];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_3 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[3];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_4 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[4];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_5 = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0[5];
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[0] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[1] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1 && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[2] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2 && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_1));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[3] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_3 && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_2));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[4] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_4 && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_3));
    _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[5] = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_5 && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_4));
  end

  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_1 = ({Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1,Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0} != 2'b00);
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_2 = ({Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2,{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1,Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0}} != 3'b000);
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_3 = ({Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_3,{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2,{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1,Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0}}} != 4'b0000);
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_range_0_to_4 = ({Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_4,{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_3,{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_2,{Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_1,Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hits_bools_0}}}} != 5'h00);
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh;
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[0];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[1];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[2];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[3];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[4];
  assign _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh[5];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_6[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException[0];
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated = ((((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated : _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_2) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_1 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_3 : _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_5)) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_2 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_6 : _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_8) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_3 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_9 : _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_11))) | ((_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_4 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_12 : 32'h00000000) | (_zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute_5 ? _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated_13 : 32'h00000000)));
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault = _zz_Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault[0];
  always @(*) begin
    Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup = (MmuPlugin_logic_satp_mode == 1'b1);
    if(when_MmuPlugin_l297) begin
      Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
    if(when_MmuPlugin_l298) begin
      if(when_MmuPlugin_l300) begin
        Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
      end
    end
  end

  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_needRefill = ((Lsu2Plugin_logic_sharedPip_stages_1_valid && (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hit)) && Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup);
  assign Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_askRefill = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_needRefill && Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded);
  assign when_MmuPlugin_l297 = ((! MmuPlugin_logic_status_mprv) && (PrivilegedPlugin_setup_privilege == 2'b11));
  assign when_MmuPlugin_l298 = (PrivilegedPlugin_setup_privilege == 2'b11);
  assign when_MmuPlugin_l300 = ((! MmuPlugin_logic_status_mprv) || (PrivilegedPlugin_logic_machine_mstatus_mpp == 2'b11));
  always @(*) begin
    PrivilegedPlugin_setup_ramWrite_valid = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_ramWrite_address = 5'bxxxxx;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_address = _zz_PrivilegedPlugin_setup_ramWrite_address;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_address = _zz_PrivilegedPlugin_setup_ramWrite_address_1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_ramWrite_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_data = _zz_PrivilegedPlugin_setup_ramWrite_data;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        PrivilegedPlugin_setup_ramWrite_data = _zz_PrivilegedPlugin_setup_ramWrite_data_1;
        if(PrivilegedPlugin_logic_decoderInterrupt_raised) begin
          PrivilegedPlugin_setup_ramWrite_data = 32'h00000000;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_ramRead_valid = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        PrivilegedPlugin_setup_ramRead_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        PrivilegedPlugin_setup_ramRead_valid = 1'b1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_setup_ramRead_address = 5'bxxxxx;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        PrivilegedPlugin_setup_ramRead_address = _zz_PrivilegedPlugin_setup_ramRead_address;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        PrivilegedPlugin_setup_ramRead_address = _zz_PrivilegedPlugin_setup_ramRead_address_1;
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_logic_interrupt_valid = 1'b0;
    if(when_PrivilegedPlugin_l631_1) begin
      if(when_PrivilegedPlugin_l637) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l637_1) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l637_2) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
    end
    if(when_PrivilegedPlugin_l631) begin
      if(when_PrivilegedPlugin_l637_3) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l637_4) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l637_5) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l637_6) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l637_7) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
      if(when_PrivilegedPlugin_l637_8) begin
        PrivilegedPlugin_logic_interrupt_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_interrupt_code = 4'bxxxx;
    if(when_PrivilegedPlugin_l631_1) begin
      if(when_PrivilegedPlugin_l637) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0001;
      end
      if(when_PrivilegedPlugin_l637_1) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0101;
      end
      if(when_PrivilegedPlugin_l637_2) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b1001;
      end
    end
    if(when_PrivilegedPlugin_l631) begin
      if(when_PrivilegedPlugin_l637_3) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0111;
      end
      if(when_PrivilegedPlugin_l637_4) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0011;
      end
      if(when_PrivilegedPlugin_l637_5) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b1011;
      end
      if(when_PrivilegedPlugin_l637_6) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0001;
      end
      if(when_PrivilegedPlugin_l637_7) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b0101;
      end
      if(when_PrivilegedPlugin_l637_8) begin
        PrivilegedPlugin_logic_interrupt_code = 4'b1001;
      end
    end
  end

  always @(*) begin
    PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'bxx;
    if(when_PrivilegedPlugin_l631_1) begin
      if(when_PrivilegedPlugin_l637) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b01;
      end
      if(when_PrivilegedPlugin_l637_1) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b01;
      end
      if(when_PrivilegedPlugin_l637_2) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b01;
      end
    end
    if(when_PrivilegedPlugin_l631) begin
      if(when_PrivilegedPlugin_l637_3) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l637_4) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l637_5) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l637_6) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l637_7) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
      if(when_PrivilegedPlugin_l637_8) begin
        PrivilegedPlugin_logic_interrupt_targetPrivilege = 2'b11;
      end
    end
  end

  assign when_PrivilegedPlugin_l631 = (PrivilegedPlugin_logic_machine_mstatus_mie || (! PrivilegedPlugin_setup_withMachinePrivilege));
  assign when_PrivilegedPlugin_l631_1 = ((PrivilegedPlugin_logic_supervisor_sstatus_sie && (! PrivilegedPlugin_setup_withMachinePrivilege)) || (! PrivilegedPlugin_setup_withSupervisorPrivilege));
  assign when_PrivilegedPlugin_l637 = ((_zz_when_PrivilegedPlugin_l637 && (1'b1 && PrivilegedPlugin_logic_machine_mideleg_ss)) && (! 1'b0));
  assign when_PrivilegedPlugin_l637_1 = ((_zz_when_PrivilegedPlugin_l637_1 && (1'b1 && PrivilegedPlugin_logic_machine_mideleg_st)) && (! 1'b0));
  assign when_PrivilegedPlugin_l637_2 = ((_zz_when_PrivilegedPlugin_l637_2 && (1'b1 && PrivilegedPlugin_logic_machine_mideleg_se)) && (! 1'b0));
  assign when_PrivilegedPlugin_l637_3 = (((PrivilegedPlugin_logic_machine_mip_mtip && PrivilegedPlugin_logic_machine_mie_mtie) && 1'b1) && (! 1'b0));
  assign when_PrivilegedPlugin_l637_4 = (((PrivilegedPlugin_logic_machine_mip_msip && PrivilegedPlugin_logic_machine_mie_msie) && 1'b1) && (! 1'b0));
  assign when_PrivilegedPlugin_l637_5 = (((PrivilegedPlugin_logic_machine_mip_meip && PrivilegedPlugin_logic_machine_mie_meie) && 1'b1) && (! 1'b0));
  assign when_PrivilegedPlugin_l637_6 = ((_zz_when_PrivilegedPlugin_l637 && 1'b1) && (! (PrivilegedPlugin_logic_machine_mideleg_ss != 1'b0)));
  assign when_PrivilegedPlugin_l637_7 = ((_zz_when_PrivilegedPlugin_l637_1 && 1'b1) && (! (PrivilegedPlugin_logic_machine_mideleg_st != 1'b0)));
  assign when_PrivilegedPlugin_l637_8 = ((_zz_when_PrivilegedPlugin_l637_2 && 1'b1) && (! (PrivilegedPlugin_logic_machine_mideleg_se != 1'b0)));
  assign PrivilegedPlugin_logic_decoderInterrupt_doIt = PrivilegedPlugin_logic_decoderInterrupt_counter[2];
  assign when_PrivilegedPlugin_l668 = (((! PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt) || (! DecoderPlugin_setup_trapReady)) || PrivilegedPlugin_logic_decoderInterrupt_raised);
  assign when_PrivilegedPlugin_l672 = (PrivilegedPlugin_logic_decoderInterrupt_doIt && (! PrivilegedPlugin_logic_decoderInterrupt_raised));
  assign PrivilegedPlugin_logic_decoderInterrupt_buffer_sample = (PrivilegedPlugin_logic_interrupt_valid && (! PrivilegedPlugin_logic_decoderInterrupt_raised));
  always @(*) begin
    PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b11;
    case(PrivilegedPlugin_logic_exception_code)
      4'b0000 : begin
        if(when_PrivilegedPlugin_l702) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b0011 : begin
        if(when_PrivilegedPlugin_l702_1) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1000 : begin
        if(when_PrivilegedPlugin_l702_2) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1001 : begin
        if(when_PrivilegedPlugin_l702_3) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1100 : begin
        if(when_PrivilegedPlugin_l702_4) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1101 : begin
        if(when_PrivilegedPlugin_l702_5) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1111 : begin
        if(when_PrivilegedPlugin_l702_6) begin
          PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_logic_exception_code = PrivilegedPlugin_logic_reschedule_payload_cause;
    if(when_PrivilegedPlugin_l689) begin
      PrivilegedPlugin_logic_exception_code[1 : 0] = PrivilegedPlugin_setup_privilege;
    end
  end

  assign when_PrivilegedPlugin_l689 = (PrivilegedPlugin_logic_reschedule_payload_cause == 4'b1011);
  assign when_PrivilegedPlugin_l702 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_iam) && (! 1'b0));
  assign when_PrivilegedPlugin_l702_1 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_bp) && (! 1'b0));
  assign when_PrivilegedPlugin_l702_2 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_eu) && (! 1'b0));
  assign when_PrivilegedPlugin_l702_3 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_es) && (! 1'b0));
  assign when_PrivilegedPlugin_l702_4 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_ipf) && (! 1'b0));
  assign when_PrivilegedPlugin_l702_5 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_lpf) && (! 1'b0));
  assign when_PrivilegedPlugin_l702_6 = ((1'b1 && PrivilegedPlugin_logic_machine_medeleg_spf) && (! 1'b0));
  assign PrivilegedPlugin_logic_exception_targetPrivilege = ((PrivilegedPlugin_setup_privilege < PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped) ? PrivilegedPlugin_logic_exception_exceptionTargetPrivilegeUncapped : PrivilegedPlugin_setup_privilege);
  assign PrivilegedPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    PrivilegedPlugin_logic_fsm_wantStart = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
        PrivilegedPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign PrivilegedPlugin_logic_fsm_wantKill = 1'b0;
  always @(*) begin
    PrivilegedPlugin_logic_fsm_trap_fire = 1'b0;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_logic_fsm_trap_fire = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_logic_fsm_xret_sourcePrivilege = PrivilegedPlugin_logic_reschedule_payload_tval[1 : 0];
  always @(*) begin
    PrivilegedPlugin_logic_fsm_xret_targetPrivilege = PrivilegedPlugin_logic_machine_mstatus_mpp;
    case(PrivilegedPlugin_logic_fsm_xret_sourcePrivilege)
      2'b01 : begin
        PrivilegedPlugin_logic_fsm_xret_targetPrivilege = {1'b0,PrivilegedPlugin_logic_supervisor_sstatus_spp};
      end
      default : begin
      end
    endcase
  end

  assign FetchPlugin_stages_0_haltRequest_PrivilegedPlugin_l968 = ((! (PrivilegedPlugin_logic_fsm_stateReg == PrivilegedPlugin_logic_fsm_enumDef_IDLE)) || (CommitPlugin_logic_reschedule_valid && CommitPlugin_logic_reschedule_trap));
  assign trap_fire = PrivilegedPlugin_logic_fsm_trap_fire;
  assign trap_code = PrivilegedPlugin_logic_fsm_trap_code;
  assign trap_interrupt = PrivilegedPlugin_logic_fsm_trap_interrupt;
  assign trap_tval = PrivilegedPlugin_logic_reschedule_payload_tval;
  always @(*) begin
    PerformanceCounterPlugin_setup_readPort_valid = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
        PerformanceCounterPlugin_setup_readPort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
        PerformanceCounterPlugin_setup_readPort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_setup_readPort_address = (5'h00 | _zz_PerformanceCounterPlugin_setup_readPort_address);
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
        PerformanceCounterPlugin_setup_readPort_address[3] = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_setup_writePort_valid = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
        PerformanceCounterPlugin_setup_writePort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
        PerformanceCounterPlugin_setup_writePort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
        PerformanceCounterPlugin_setup_writePort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_setup_writePort_address = (5'h00 | _zz_PerformanceCounterPlugin_setup_writePort_address);
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
        PerformanceCounterPlugin_setup_writePort_address[3] = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
        PerformanceCounterPlugin_setup_writePort_address = (5'h00 | _zz_PerformanceCounterPlugin_setup_writePort_address_1);
        PerformanceCounterPlugin_setup_writePort_address[3] = PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_high;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_setup_writePort_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
        PerformanceCounterPlugin_setup_writePort_data = _zz_PerformanceCounterPlugin_setup_writePort_data[31:0];
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
        PerformanceCounterPlugin_setup_writePort_data = _zz_PerformanceCounterPlugin_setup_writePort_data_1;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
        PerformanceCounterPlugin_setup_writePort_data = EU0_CsrAccessPlugin_setup_onWriteBits;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_fsm_calc = {_zz_PerformanceCounterPlugin_logic_fsm_calc,_zz_PerformanceCounterPlugin_logic_fsm_calc_3};
  assign PerformanceCounterPlugin_logic_flusher_hits = {_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6[5],{_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5[5],{_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4[5],{_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3[5],{_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2[5],{_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_1[5],_zz_PerformanceCounterPlugin_logic_fsm_counterReaded[5]}}}}}};
  assign PerformanceCounterPlugin_logic_flusher_hit = (|PerformanceCounterPlugin_logic_flusher_hits);
  assign PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input = PerformanceCounterPlugin_logic_flusher_hits;
  assign PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked = (PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input & (~ _zz_PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked));
  assign PerformanceCounterPlugin_logic_flusher_oh = PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked;
  assign _zz_PerformanceCounterPlugin_logic_flusher_sel = PerformanceCounterPlugin_logic_flusher_oh[3];
  assign _zz_PerformanceCounterPlugin_logic_flusher_sel_1 = PerformanceCounterPlugin_logic_flusher_oh[5];
  assign _zz_PerformanceCounterPlugin_logic_flusher_sel_2 = PerformanceCounterPlugin_logic_flusher_oh[6];
  assign _zz_PerformanceCounterPlugin_logic_flusher_sel_3 = ((PerformanceCounterPlugin_logic_flusher_oh[1] || _zz_PerformanceCounterPlugin_logic_flusher_sel) || _zz_PerformanceCounterPlugin_logic_flusher_sel_1);
  assign _zz_PerformanceCounterPlugin_logic_flusher_sel_4 = ((PerformanceCounterPlugin_logic_flusher_oh[2] || _zz_PerformanceCounterPlugin_logic_flusher_sel) || _zz_PerformanceCounterPlugin_logic_flusher_sel_2);
  assign _zz_PerformanceCounterPlugin_logic_flusher_sel_5 = ((PerformanceCounterPlugin_logic_flusher_oh[4] || _zz_PerformanceCounterPlugin_logic_flusher_sel_1) || _zz_PerformanceCounterPlugin_logic_flusher_sel_2);
  assign PerformanceCounterPlugin_logic_flusher_sel = {_zz_PerformanceCounterPlugin_logic_flusher_sel_5,{_zz_PerformanceCounterPlugin_logic_flusher_sel_4,_zz_PerformanceCounterPlugin_logic_flusher_sel_3}};
  assign PerformanceCounterPlugin_logic_fsm_flusherCmd_valid = PerformanceCounterPlugin_logic_flusher_hit;
  assign PerformanceCounterPlugin_logic_fsm_flusherCmd_payload_address = PerformanceCounterPlugin_logic_flusher_sel;
  assign PerformanceCounterPlugin_logic_fsm_csrReadCmd_fire = (PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid && PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready);
  always @(*) begin
    PerformanceCounterPlugin_logic_csrRead_requested = 1'b0;
    if(when_CsrAccessPlugin_l244) begin
      PerformanceCounterPlugin_logic_csrRead_requested = 1'b1;
    end
  end

  assign PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid = (PerformanceCounterPlugin_logic_csrRead_requested && (! PerformanceCounterPlugin_logic_csrRead_fired));
  assign PerformanceCounterPlugin_logic_fsm_csrReadCmd_payload_address = EU0_CsrAccessPlugin_setup_onReadAddress[2 : 0];
  assign when_PerformanceCounterPlugin_l253 = ((! PerformanceCounterPlugin_logic_csrRead_fired) || (! PerformanceCounterPlugin_logic_fsm_done));
  assign PerformanceCounterPlugin_logic_fsm_csrWriteCmd_fire = (PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid && PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready);
  assign PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address = EU0_CsrAccessPlugin_setup_onWriteAddress[2 : 0];
  assign PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_high = EU0_CsrAccessPlugin_setup_onWriteAddress[7];
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid = 1'b0;
    if(when_CsrAccessPlugin_l325) begin
      if(when_PerformanceCounterPlugin_l273) begin
        PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid = 1'b1;
      end
    end
  end

  assign when_PerformanceCounterPlugin_l268 = (EU0_CsrAccessPlugin_setup_onDecodeWrite && ((EU0_CsrAccessPlugin_setup_onDecodeAddress & 12'hf60) == 12'hc00));
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_IO = (Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED[31 : 28] == 4'b0001);
  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO = (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_hit);
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO = 1'b0;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineTranslated;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED = Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_EXECUTE = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute && (! (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser && (PrivilegedPlugin_setup_privilege == 2'b01))));
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_EXECUTE = 1'b1;
    end
    if(when_MmuPlugin_l326) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_EXECUTE = 1'b0;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ = (Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ = 1'b1;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_WRITE = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_WRITE = 1'b1;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT = ((Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineException || ((Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser && (PrivilegedPlugin_setup_privilege == 2'b01)) && (! MmuPlugin_logic_status_sum))) || ((! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAllowUser) && (PrivilegedPlugin_setup_privilege == 2'b00)));
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT = 1'b0;
    end
  end

  always @(*) begin
    if(Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup) begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_lineAccessFault;
    end else begin
      Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT = 1'b0;
    end
  end

  assign when_MmuPlugin_l326 = (! (Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED[31 : 28] != 4'b0001));
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_BYPASS_TRANSLATION = (! Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_requireMmuLockup);
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_OH = Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_oh;
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_0 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_1 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_2 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_3 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[11 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_4 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[21 : 0]};
  assign Lsu2Plugin_logic_sharedPip_stages_1_MMU_WAYS_PHYSICAL_5 = {Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_physicalAddress,Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION[21 : 0]};
  assign FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL = 1'b1;
  assign FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded = ((FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL && (! FetchCachePlugin_setup_translationStorage_logic_refillOngoing)) && FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg);
  assign when_MmuPlugin_l260_2 = (FetchPlugin_stages_1_isRemoved || (! (FetchPlugin_stages_1_valid && (! FetchPlugin_stages_1_ready))));
  assign FetchCachePlugin_logic_translationPort_logic_read_0_readAddress = FetchPlugin_stages_1_Fetch_FETCH_PC[16 : 12];
  assign _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid = _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_0_port1;
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[0];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_pageFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[1];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_accessFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[2];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[17 : 3];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[37 : 18];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowRead = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[38];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowWrite = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[39];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowExecute = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[40];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_0_allowUser = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid[41];
  always @(*) begin
    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[0] = (FetchPlugin_stages_1_MMU_L0_ENTRIES_0_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 17]);
    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[1] = (FetchPlugin_stages_1_MMU_L0_ENTRIES_1_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 17]);
    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[2] = (FetchPlugin_stages_1_MMU_L0_ENTRIES_2_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 17]);
    FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[3] = (FetchPlugin_stages_1_MMU_L0_ENTRIES_3_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 17]);
  end

  always @(*) begin
    FetchPlugin_stages_1_MMU_L0_HITS[0] = (FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[0] && FetchPlugin_stages_1_MMU_L0_ENTRIES_0_valid);
    FetchPlugin_stages_1_MMU_L0_HITS[1] = (FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[1] && FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid);
    FetchPlugin_stages_1_MMU_L0_HITS[2] = (FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[2] && FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid);
    FetchPlugin_stages_1_MMU_L0_HITS[3] = (FetchPlugin_stages_1_MMU_L0_HITS_PRE_VALID[3] && FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid);
  end

  assign _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid = _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_1_port1;
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[0];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_pageFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[1];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_accessFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[2];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[17 : 3];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[37 : 18];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowRead = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[38];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowWrite = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[39];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowExecute = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[40];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_1_allowUser = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_1_valid[41];
  assign _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid = _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_2_port1;
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[0];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_pageFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[1];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_accessFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[2];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[17 : 3];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[37 : 18];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowRead = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[38];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowWrite = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[39];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowExecute = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[40];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_2_allowUser = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_2_valid[41];
  assign _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid = _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_ways_3_port1;
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[0];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_pageFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[1];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_accessFault = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[2];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[17 : 3];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[37 : 18];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowRead = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[38];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowWrite = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[39];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowExecute = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[40];
  assign FetchPlugin_stages_1_MMU_L0_ENTRIES_3_allowUser = _zz_FetchPlugin_stages_1_MMU_L0_ENTRIES_3_valid[41];
  assign FetchCachePlugin_logic_translationPort_logic_read_1_readAddress = FetchPlugin_stages_1_Fetch_FETCH_PC[26 : 22];
  assign _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid = _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_0_port1;
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[0];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_pageFault = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[1];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_accessFault = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[2];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[7 : 3];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[17 : 8];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowRead = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[18];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowWrite = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[19];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowExecute = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[20];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_0_allowUser = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid[21];
  always @(*) begin
    FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID[0] = (FetchPlugin_stages_1_MMU_L1_ENTRIES_0_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 27]);
    FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID[1] = (FetchPlugin_stages_1_MMU_L1_ENTRIES_1_virtualAddress == FetchPlugin_stages_1_Fetch_FETCH_PC[31 : 27]);
  end

  always @(*) begin
    FetchPlugin_stages_1_MMU_L1_HITS[0] = (FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID[0] && FetchPlugin_stages_1_MMU_L1_ENTRIES_0_valid);
    FetchPlugin_stages_1_MMU_L1_HITS[1] = (FetchPlugin_stages_1_MMU_L1_HITS_PRE_VALID[1] && FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid);
  end

  assign _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid = _zz_FetchCachePlugin_setup_translationStorage_logic_sl_1_ways_1_port1;
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[0];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_pageFault = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[1];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_accessFault = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[2];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_virtualAddress = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[7 : 3];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_physicalAddress = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[17 : 8];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowRead = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[18];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowWrite = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[19];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowExecute = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[20];
  assign FetchPlugin_stages_1_MMU_L1_ENTRIES_1_allowUser = _zz_FetchPlugin_stages_1_MMU_L1_ENTRIES_1_valid[21];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits = {FetchPlugin_stages_1_MMU_L1_HITS,FetchPlugin_stages_1_MMU_L0_HITS};
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hit = (|FetchCachePlugin_logic_translationPort_logic_ctrl_hits);
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0 = FetchCachePlugin_logic_translationPort_logic_ctrl_hits;
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[1];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[2];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_3 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[3];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_4 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[4];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_5 = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0[5];
  always @(*) begin
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[0] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[1] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1 && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[2] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2 && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_1));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[3] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_3 && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_2));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[4] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_4 && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_3));
    _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh[5] = (FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_5 && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_4));
  end

  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_1 = ({FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0} != 2'b00);
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_2 = ({FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2,{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0}} != 3'b000);
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_3 = ({FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_3,{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2,{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0}}} != 4'b0000);
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_hits_range_0_to_4 = ({FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_4,{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_3,{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_2,{FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchCachePlugin_logic_translationPort_logic_ctrl_hits_bools_0}}}} != 5'h00);
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_oh = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_oh;
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[0];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[1];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[2];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[3];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[4];
  assign _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 = FetchCachePlugin_logic_translationPort_logic_ctrl_oh[5];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_6[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineException = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineException[0];
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated = ((((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated : _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_2) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_3 : _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_5)) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_6 : _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_8) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_9 : _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_11))) | ((_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_4 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_12 : 32'h00000000) | (_zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute_5 ? _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated_13 : 32'h00000000)));
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault = _zz_FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault[0];
  always @(*) begin
    FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup = (MmuPlugin_logic_satp_mode == 1'b1);
    if(when_MmuPlugin_l297_1) begin
      FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
    if(when_MmuPlugin_l298_1) begin
      FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
  end

  assign FetchCachePlugin_logic_translationPort_logic_ctrl_needRefill = ((FetchPlugin_stages_1_valid && (! FetchCachePlugin_logic_translationPort_logic_ctrl_hit)) && FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup);
  assign FetchCachePlugin_logic_translationPort_logic_ctrl_askRefill = (FetchCachePlugin_logic_translationPort_logic_ctrl_needRefill && FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded);
  assign when_MmuPlugin_l297_1 = ((! MmuPlugin_logic_status_mprv) && (PrivilegedPlugin_setup_privilege == 2'b11));
  assign when_MmuPlugin_l298_1 = (PrivilegedPlugin_setup_privilege == 2'b11);
  assign FetchPlugin_stages_1_MMU_IO = (FetchPlugin_stages_1_MMU_TRANSLATED[31 : 28] == 4'b0001);
  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_REDO = (! FetchCachePlugin_logic_translationPort_logic_ctrl_hit);
    end else begin
      FetchPlugin_stages_1_MMU_REDO = 1'b0;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_TRANSLATED = FetchCachePlugin_logic_translationPort_logic_ctrl_lineTranslated;
    end else begin
      FetchPlugin_stages_1_MMU_TRANSLATED = FetchPlugin_stages_1_Fetch_FETCH_PC;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_ALLOW_EXECUTE = (FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute && (! (FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser && (PrivilegedPlugin_setup_privilege == 2'b01))));
    end else begin
      FetchPlugin_stages_1_MMU_ALLOW_EXECUTE = 1'b1;
    end
    if(when_MmuPlugin_l326_1) begin
      FetchPlugin_stages_1_MMU_ALLOW_EXECUTE = 1'b0;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_ALLOW_READ = (FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      FetchPlugin_stages_1_MMU_ALLOW_READ = 1'b1;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_ALLOW_WRITE = FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      FetchPlugin_stages_1_MMU_ALLOW_WRITE = 1'b1;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_PAGE_FAULT = ((FetchCachePlugin_logic_translationPort_logic_ctrl_lineException || ((FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser && (PrivilegedPlugin_setup_privilege == 2'b01)) && (! MmuPlugin_logic_status_sum))) || ((! FetchCachePlugin_logic_translationPort_logic_ctrl_lineAllowUser) && (PrivilegedPlugin_setup_privilege == 2'b00)));
    end else begin
      FetchPlugin_stages_1_MMU_PAGE_FAULT = 1'b0;
    end
  end

  always @(*) begin
    if(FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      FetchPlugin_stages_1_MMU_ACCESS_FAULT = FetchCachePlugin_logic_translationPort_logic_ctrl_lineAccessFault;
    end else begin
      FetchPlugin_stages_1_MMU_ACCESS_FAULT = 1'b0;
    end
  end

  assign when_MmuPlugin_l326_1 = (! (FetchPlugin_stages_1_MMU_TRANSLATED[31 : 28] != 4'b0001));
  assign FetchPlugin_stages_1_MMU_BYPASS_TRANSLATION = (! FetchCachePlugin_logic_translationPort_logic_ctrl_requireMmuLockup);
  assign FetchPlugin_stages_1_MMU_WAYS_OH = FetchCachePlugin_logic_translationPort_logic_ctrl_oh;
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_0 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_0_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_1 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_1_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_2 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_2_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_3 = {FetchPlugin_stages_1_MMU_L0_ENTRIES_3_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[11 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_4 = {FetchPlugin_stages_1_MMU_L1_ENTRIES_0_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[21 : 0]};
  assign FetchPlugin_stages_1_MMU_WAYS_PHYSICAL_5 = {FetchPlugin_stages_1_MMU_L1_ENTRIES_1_physicalAddress,FetchPlugin_stages_1_Fetch_FETCH_PC[21 : 0]};
  assign MmuPlugin_logic_refill_wantExit = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_wantStart = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
        MmuPlugin_logic_refill_wantStart = 1'b1;
      end
    endcase
  end

  assign MmuPlugin_logic_refill_wantKill = 1'b0;
  assign MmuPlugin_logic_refill_busy = (! (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_enumDef_IDLE));
  assign _zz_Lsu2Plugin_setup_translationStorage_logic_sl_0_write_mask = MmuPlugin_logic_refill_portOhReg[0];
  assign _zz_FetchCachePlugin_setup_translationStorage_logic_sl_0_write_mask = MmuPlugin_logic_refill_portOhReg[1];
  assign MmuPlugin_logic_refill_portsRequests = {FetchCachePlugin_logic_translationPort_logic_ctrl_askRefill,Lsu2Plugin_logic_sharedPip_translationPort_logic_ctrl_askRefill};
  always @(*) begin
    MmuPlugin_logic_refill_portsRequest = (|MmuPlugin_logic_refill_portsRequests);
    if(when_MmuPlugin_l492) begin
      MmuPlugin_logic_refill_portsRequest = 1'b0;
    end
    if(when_MmuPlugin_l505) begin
      MmuPlugin_logic_refill_portsRequest = 1'b0;
    end
  end

  assign MmuPlugin_logic_refill_portsRequests_ohFirst_input = MmuPlugin_logic_refill_portsRequests;
  assign MmuPlugin_logic_refill_portsRequests_ohFirst_masked = (MmuPlugin_logic_refill_portsRequests_ohFirst_input & (~ _zz_MmuPlugin_logic_refill_portsRequests_ohFirst_masked));
  assign MmuPlugin_logic_refill_portsOh = MmuPlugin_logic_refill_portsRequests_ohFirst_masked;
  assign MmuPlugin_logic_refill_portsAddress = ((MmuPlugin_logic_refill_portsOh_regNext[0] ? _zz_MmuPlugin_logic_refill_portsAddress : 32'h00000000) | (MmuPlugin_logic_refill_portsOh_regNext[1] ? _zz_MmuPlugin_logic_refill_portsAddress_1 : 32'h00000000));
  always @(*) begin
    MmuPlugin_logic_refill_cacheRefillSet = 2'b00;
    if(when_MmuPlugin_l388) begin
      MmuPlugin_logic_refill_cacheRefillSet = MmuPlugin_setup_cacheLoad_rsp_payload_refillSlot;
    end
  end

  always @(*) begin
    MmuPlugin_logic_refill_cacheRefillAnySet = 1'b0;
    if(when_MmuPlugin_l388) begin
      MmuPlugin_logic_refill_cacheRefillAnySet = MmuPlugin_setup_cacheLoad_rsp_payload_refillSlotAny;
    end
  end

  assign FetchCachePlugin_logic_translationPort_wake = MmuPlugin_logic_refill_doWake;
  assign Lsu2Plugin_logic_sharedPip_translationPort_wake = MmuPlugin_logic_refill_doWake;
  assign MmuPlugin_logic_refill_load_readed = MmuPlugin_logic_refill_load_rsp_payload_data[31 : 0];
  assign when_MmuPlugin_l388 = (MmuPlugin_setup_cacheLoad_rsp_valid && MmuPlugin_setup_cacheLoad_rsp_payload_redo);
  always @(*) begin
    MmuPlugin_setup_cacheLoad_cmd_valid = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
        if(when_MmuPlugin_l452) begin
          MmuPlugin_setup_cacheLoad_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
        if(when_MmuPlugin_l452_1) begin
          MmuPlugin_setup_cacheLoad_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_setup_cacheLoad_cmd_payload_virtual = MmuPlugin_logic_refill_load_address;
  assign MmuPlugin_setup_cacheLoad_cmd_payload_size = 2'b10;
  assign MmuPlugin_setup_cacheLoad_cmd_payload_redoOnDataHazard = 1'b1;
  assign MmuPlugin_setup_cacheLoad_cmd_payload_unlocked = 1'b0;
  assign MmuPlugin_setup_cacheLoad_cmd_payload_unique = 1'b0;
  assign MmuPlugin_setup_cacheLoad_translated_physical = MmuPlugin_logic_refill_load_address;
  assign MmuPlugin_setup_cacheLoad_translated_abord = 1'b0;
  assign MmuPlugin_setup_cacheLoad_cancels = 3'b000;
  assign _zz_MmuPlugin_logic_refill_load_flags_V = MmuPlugin_logic_refill_load_readed;
  assign MmuPlugin_logic_refill_load_flags_V = _zz_MmuPlugin_logic_refill_load_flags_V[0];
  assign MmuPlugin_logic_refill_load_flags_R = _zz_MmuPlugin_logic_refill_load_flags_V[1];
  assign MmuPlugin_logic_refill_load_flags_W = _zz_MmuPlugin_logic_refill_load_flags_V[2];
  assign MmuPlugin_logic_refill_load_flags_X = _zz_MmuPlugin_logic_refill_load_flags_V[3];
  assign MmuPlugin_logic_refill_load_flags_U = _zz_MmuPlugin_logic_refill_load_flags_V[4];
  assign MmuPlugin_logic_refill_load_flags_G = _zz_MmuPlugin_logic_refill_load_flags_V[5];
  assign MmuPlugin_logic_refill_load_flags_A = _zz_MmuPlugin_logic_refill_load_flags_V[6];
  assign MmuPlugin_logic_refill_load_flags_D = _zz_MmuPlugin_logic_refill_load_flags_V[7];
  assign MmuPlugin_logic_refill_load_leaf = (MmuPlugin_logic_refill_load_flags_R || MmuPlugin_logic_refill_load_flags_X);
  always @(*) begin
    MmuPlugin_logic_refill_load_exception = ((((! MmuPlugin_logic_refill_load_flags_V) || ((! MmuPlugin_logic_refill_load_flags_R) && MmuPlugin_logic_refill_load_flags_W)) || MmuPlugin_logic_refill_load_rsp_payload_fault) || ((! MmuPlugin_logic_refill_load_leaf) && ((MmuPlugin_logic_refill_load_flags_D || MmuPlugin_logic_refill_load_flags_A) || MmuPlugin_logic_refill_load_flags_U)));
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(when_MmuPlugin_l461) begin
          MmuPlugin_logic_refill_load_exception = 1'b1;
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_load_levelException_0 = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_load_levelException_1 = 1'b0;
    if(when_MmuPlugin_l416) begin
      MmuPlugin_logic_refill_load_levelException_1 = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_nextLevelBase = 32'h00000000;
    MmuPlugin_logic_refill_load_nextLevelBase[21 : 12] = MmuPlugin_logic_refill_load_readed[19 : 10];
    MmuPlugin_logic_refill_load_nextLevelBase[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 = 32'h00000000;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[21 : 12] = MmuPlugin_logic_refill_load_readed[19 : 10];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 = 32'h00000000;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[21 : 12] = MmuPlugin_logic_refill_virtual[21 : 12];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  assign when_MmuPlugin_l416 = (MmuPlugin_logic_refill_load_readed[19 : 10] != 10'h000);
  always @(*) begin
    MmuPlugin_logic_invalidate_canStart = 1'b1;
    if(when_MmuPlugin_l511) begin
      MmuPlugin_logic_invalidate_canStart = 1'b0;
    end
  end

  assign MmuPlugin_logic_invalidate_done = MmuPlugin_logic_invalidate_counter[5];
  assign when_MmuPlugin_l492 = (! MmuPlugin_logic_invalidate_done);
  assign FetchPlugin_stages_0_haltRequest_MmuPlugin_l503 = ((! MmuPlugin_logic_invalidate_done) || MmuPlugin_logic_invalidate_requested);
  assign when_MmuPlugin_l505 = (MmuPlugin_logic_invalidate_requested && MmuPlugin_logic_invalidate_canStart);
  assign when_MmuPlugin_l511 = (MmuPlugin_logic_refill_busy || (Lsu2Plugin_setup_postCommitBusy != 1'b0));
  assign when_MmuPlugin_l515 = (MmuPlugin_logic_invalidate_done && (! MmuPlugin_logic_invalidate_done_regNext));
  assign EU0_CsrAccessPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_wantStart = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
        EU0_CsrAccessPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign EU0_CsrAccessPlugin_logic_fsm_wantKill = 1'b0;
  assign Lsu2Plugin_logic_sharedPip_stages_3_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_2_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_1_isRemoved = (Lsu2Plugin_logic_sharedPip_stages_1_isFlushed || Lsu2Plugin_logic_sharedPip_stages_1_isThrown);
  assign Lsu2Plugin_logic_sharedPip_stages_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_1_isThrown = 1'b0;
  assign Lsu2Plugin_logic_sharedPip_stages_0_isRemoved = (Lsu2Plugin_logic_sharedPip_stages_0_isFlushed || Lsu2Plugin_logic_sharedPip_stages_0_isThrown);
  assign Lsu2Plugin_logic_sharedPip_stages_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_0_isThrown = 1'b0;
  always @(*) begin
    _zz_Lsu2Plugin_logic_sharedPip_stages_1_valid = Lsu2Plugin_logic_sharedPip_stages_0_valid;
    if(when_Pipeline_l278) begin
      _zz_Lsu2Plugin_logic_sharedPip_stages_1_valid = 1'b0;
    end
  end

  always @(*) begin
    Lsu2Plugin_logic_sharedPip_stages_0_ready = 1'b1;
    if(when_Pipeline_l278) begin
      Lsu2Plugin_logic_sharedPip_stages_0_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278 = (Lsu2Plugin_logic_sharedPip_stages_0_haltRequest_Lsu2Plugin_l990 != 1'b0);
  assign Lsu2Plugin_logic_sharedPip_stages_1_ready = 1'b1;
  assign Lsu2Plugin_logic_sharedPip_stages_2_ready = 1'b1;
  assign Lsu2Plugin_logic_sharedPip_stages_3_ready = 1'b1;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_valid = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_valid;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_data = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_data;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_fault = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_fault;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_redo = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_redo;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlot = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlot;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_resulting_payload_refillSlotAny = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny;
  assign Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_resulting = Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
  assign Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_resulting = Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED_overloaded;
  assign Lsu2Plugin_logic_lqSqArbitration_s1_isRemoved = (Lsu2Plugin_logic_lqSqArbitration_s1_isFlushed || Lsu2Plugin_logic_lqSqArbitration_s1_isThrown);
  assign Lsu2Plugin_logic_lqSqArbitration_s1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_lqSqArbitration_s1_isThrown = 1'b0;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign Lsu2Plugin_logic_lqSqArbitration_s0_ready = Lsu2Plugin_logic_lqSqArbitration_s0_ready_output;
  always @(*) begin
    Lsu2Plugin_logic_lqSqArbitration_s1_ready = 1'b1;
    if(when_Pipeline_l278_1) begin
      Lsu2Plugin_logic_lqSqArbitration_s1_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_1 = ({Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l842,Lsu2Plugin_logic_lqSqArbitration_s1_haltRequest_Lsu2Plugin_l834} != 2'b00);
  always @(*) begin
    Lsu2Plugin_logic_lqSqArbitration_s0_ready_output = Lsu2Plugin_logic_lqSqArbitration_s1_ready;
    if(when_Connection_l74) begin
      Lsu2Plugin_logic_lqSqArbitration_s0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74 = (! Lsu2Plugin_logic_lqSqArbitration_s1_valid);
  always @(*) begin
    Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_stateReg;
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
        if(when_Lsu2Plugin_l1704) begin
          if(when_Lsu2Plugin_l1705) begin
            Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY;
          end
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
        if(Lsu2Plugin_setup_cacheLoad_cmd_fire) begin
          Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP;
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
        if(Lsu2Plugin_setup_cacheLoad_rsp_valid) begin
          if(Lsu2Plugin_setup_cacheLoad_rsp_payload_redo) begin
            Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD;
          end else begin
            if(Lsu2Plugin_setup_cacheLoad_rsp_payload_fault) begin
              Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_TRAP;
            end else begin
              Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_ALU;
            end
          end
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
        if(when_Lsu2Plugin_l1715) begin
          if(Lsu2Plugin_logic_special_storeSc) begin
            Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_ALU;
          end else begin
            Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD;
          end
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
        Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
        Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_SYNC;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
        if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
          Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_IDLE;
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
        Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_IDLE;
      end
      default : begin
      end
    endcase
    if(Lsu2Plugin_logic_special_atomic_wantStart) begin
      Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_IDLE;
    end
    if(Lsu2Plugin_logic_special_atomic_wantKill) begin
      Lsu2Plugin_logic_special_atomic_stateNext = Lsu2Plugin_logic_special_atomic_enumDef_BOOT;
    end
  end

  assign when_Lsu2Plugin_l1704 = (Lsu2Plugin_logic_special_enabled && Lsu2Plugin_logic_special_isAtomic);
  assign when_Lsu2Plugin_l1705 = (Lsu2Plugin_logic_sq_ptr_commit == Lsu2Plugin_logic_sq_ptr_free);
  assign Lsu2Plugin_setup_cacheLoad_cmd_fire = (Lsu2Plugin_setup_cacheLoad_cmd_valid && Lsu2Plugin_setup_cacheLoad_cmd_ready);
  assign when_Lsu2Plugin_l1715 = (&Lsu2Plugin_logic_special_atomic_lockDelayCounter);
  assign when_Lsu2Plugin_l1824 = (Lsu2Plugin_logic_special_storeSc && (! Lsu2Plugin_logic_special_atomic_gotReservation));
  assign when_StateMachine_l253 = ((! ((Lsu2Plugin_logic_special_atomic_stateReg & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) != 9'b000000000)) && ((Lsu2Plugin_logic_special_atomic_stateNext & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) != 9'b000000000));
  assign when_StateMachine_l253_1 = ((! ((Lsu2Plugin_logic_special_atomic_stateReg & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) != 9'b000000000)) && ((Lsu2Plugin_logic_special_atomic_stateNext & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) != 9'b000000000));
  always @(*) begin
    MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_stateReg;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
        if(MmuPlugin_logic_refill_portsRequest) begin
          MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_INIT;
        end
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
        MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_1;
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
        if(when_MmuPlugin_l452) begin
          if(MmuPlugin_setup_cacheLoad_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_RSP_0;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
        if(when_MmuPlugin_l452_1) begin
          if(MmuPlugin_setup_cacheLoad_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_RSP_1;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_0;
          end else begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_IDLE;
          end
        end
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_1;
          end else begin
            if(when_MmuPlugin_l469) begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_IDLE;
            end else begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_CMD_0;
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(MmuPlugin_logic_refill_wantStart) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_IDLE;
    end
    if(MmuPlugin_logic_refill_wantKill) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_enumDef_BOOT;
    end
  end

  assign when_MmuPlugin_l452 = ((MmuPlugin_logic_refill_cacheRefill == 2'b00) && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l452_1 = ((MmuPlugin_logic_refill_cacheRefill == 2'b00) && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l461 = (! MmuPlugin_logic_refill_load_leaf);
  assign when_MmuPlugin_l469 = (MmuPlugin_logic_refill_load_leaf || MmuPlugin_logic_refill_load_exception);
  assign MmuPlugin_logic_refill_doWake = (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_enumDef_IDLE);
  assign CsrRamPlugin_logic_flush_done = CsrRamPlugin_logic_flush_counter[5];
  assign CsrRamPlugin_setup_initPort_valid = (! CsrRamPlugin_logic_flush_done);
  assign CsrRamPlugin_setup_initPort_address = CsrRamPlugin_logic_flush_counter[4:0];
  assign CsrRamPlugin_setup_initPort_data = 32'h00000000;
  assign when_CsrRamPlugin_l61 = ((! CsrRamPlugin_logic_flush_done) && CsrRamPlugin_setup_initPort_ready);
  assign CsrRamPlugin_logic_writeLogic_hits = {CsrRamPlugin_setup_initPort_valid,{PrivilegedPlugin_setup_ramWrite_valid,{PerformanceCounterPlugin_setup_writePort_valid,EU0_CsrAccessPlugin_logic_ramWritePort_valid}}};
  assign CsrRamPlugin_logic_writeLogic_hit = (|CsrRamPlugin_logic_writeLogic_hits);
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_input = CsrRamPlugin_logic_writeLogic_hits;
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_writeLogic_oh = CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  assign _zz_PerformanceCounterPlugin_setup_writePort_ready = CsrRamPlugin_logic_writeLogic_oh[1];
  assign _zz_PrivilegedPlugin_setup_ramWrite_ready = CsrRamPlugin_logic_writeLogic_oh[2];
  assign _zz_CsrRamPlugin_setup_initPort_ready = CsrRamPlugin_logic_writeLogic_oh[3];
  assign _zz_CsrRamPlugin_logic_writeLogic_sel = (_zz_PerformanceCounterPlugin_setup_writePort_ready || _zz_CsrRamPlugin_setup_initPort_ready);
  assign _zz_CsrRamPlugin_logic_writeLogic_sel_1 = (_zz_PrivilegedPlugin_setup_ramWrite_ready || _zz_CsrRamPlugin_setup_initPort_ready);
  assign CsrRamPlugin_logic_writeLogic_sel = {_zz_CsrRamPlugin_logic_writeLogic_sel_1,_zz_CsrRamPlugin_logic_writeLogic_sel};
  assign CsrRamPlugin_logic_writeLogic_port_valid = CsrRamPlugin_logic_writeLogic_hit;
  assign CsrRamPlugin_logic_writeLogic_port_payload_address = _zz_CsrRamPlugin_logic_writeLogic_port_payload_address;
  assign CsrRamPlugin_logic_writeLogic_port_payload_data = _zz_CsrRamPlugin_logic_writeLogic_port_payload_data;
  assign EU0_CsrAccessPlugin_logic_ramWritePort_ready = CsrRamPlugin_logic_writeLogic_oh[0];
  assign PerformanceCounterPlugin_setup_writePort_ready = _zz_PerformanceCounterPlugin_setup_writePort_ready;
  assign PrivilegedPlugin_setup_ramWrite_ready = _zz_PrivilegedPlugin_setup_ramWrite_ready;
  assign CsrRamPlugin_setup_initPort_ready = _zz_CsrRamPlugin_setup_initPort_ready;
  assign CsrRamPlugin_logic_readLogic_hits = {PrivilegedPlugin_setup_ramRead_valid,{PerformanceCounterPlugin_setup_readPort_valid,EU0_CsrAccessPlugin_logic_ramReadPort_valid}};
  assign CsrRamPlugin_logic_readLogic_hit = (|CsrRamPlugin_logic_readLogic_hits);
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_input = CsrRamPlugin_logic_readLogic_hits;
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_readLogic_oh = CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  assign _zz_PerformanceCounterPlugin_setup_readPort_ready = CsrRamPlugin_logic_readLogic_oh[1];
  assign _zz_PrivilegedPlugin_setup_ramRead_ready = CsrRamPlugin_logic_readLogic_oh[2];
  assign CsrRamPlugin_logic_readLogic_sel = {_zz_PrivilegedPlugin_setup_ramRead_ready,_zz_PerformanceCounterPlugin_setup_readPort_ready};
  assign CsrRamPlugin_logic_readLogic_port_data = _zz_CsrRamPlugin_logic_mem_port1;
  assign CsrRamPlugin_logic_readLogic_port_address = _zz_CsrRamPlugin_logic_readLogic_port_address;
  assign EU0_CsrAccessPlugin_logic_ramReadPort_ready = CsrRamPlugin_logic_readLogic_oh[0];
  assign PerformanceCounterPlugin_setup_readPort_ready = _zz_PerformanceCounterPlugin_setup_readPort_ready;
  assign PrivilegedPlugin_setup_ramRead_ready = _zz_PrivilegedPlugin_setup_ramRead_ready;
  assign EU0_CsrAccessPlugin_logic_ramReadPort_data = CsrRamPlugin_logic_readLogic_port_data;
  assign PerformanceCounterPlugin_setup_readPort_data = CsrRamPlugin_logic_readLogic_port_data;
  assign PrivilegedPlugin_setup_ramRead_data = CsrRamPlugin_logic_readLogic_port_data;
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_immZero = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[19 : 15] == 5'h00);
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_srcZero = (EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_IMM ? EU0_CsrAccessPlugin_logic_fsm_startLogic_immZero : (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[19 : 15] == 5'h00));
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_csrWrite = (! (EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK && EU0_CsrAccessPlugin_logic_fsm_startLogic_srcZero));
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_csrRead = (! ((! EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK) && (! EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD)));
  assign COMB_CSR_773 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h305);
  assign COMB_CSR_835 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h343);
  assign COMB_CSR_833 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h341);
  assign COMB_CSR_832 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h340);
  assign COMB_CSR_3857 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hf11);
  assign COMB_CSR_3858 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hf12);
  assign COMB_CSR_3859 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hf13);
  assign COMB_CSR_3860 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hf14);
  assign COMB_CSR_769 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h301);
  assign COMB_CSR_834 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h342);
  assign COMB_CSR_768 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h300);
  assign COMB_CSR_836 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h344);
  assign COMB_CSR_772 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h304);
  assign COMB_CSR_770 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h302);
  assign COMB_CSR_771 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h303);
  assign COMB_CSR_261 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h105);
  assign COMB_CSR_323 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h143);
  assign COMB_CSR_321 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h141);
  assign COMB_CSR_320 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h140);
  assign COMB_CSR_322 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h142);
  assign COMB_CSR_256 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h100);
  assign COMB_CSR_260 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h104);
  assign COMB_CSR_324 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h144);
  assign COMB_CSR_262 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h106);
  assign COMB_CSR_774 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h306);
  assign COMB_CSR_ = ({(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h33f),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb9f),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hb1f),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h33e),{(_zz_COMB_CSR_ == _zz_COMB_CSR__1),{_zz_COMB_CSR__2,{_zz_COMB_CSR__3,_zz_COMB_CSR__4}}}}}}} != 87'h0000000000000000000000);
  assign COMB_CSR_803 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h323);
  assign COMB_CSR_804 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h324);
  assign COMB_CSR_805 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h325);
  assign COMB_CSR_806 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h326);
  assign COMB_CSR_384 = (EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'h180);
  assign COMB_CSR_PerformanceCounterPlugin_logic_csrFilter = ({(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc86),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc85),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc84),{(EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20] == 12'hc83),{(_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter == _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_1),{_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_2,{_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_3,_zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_4}}}}}}} != 24'h000000);
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented = ({COMB_CSR_PerformanceCounterPlugin_logic_csrFilter,{COMB_CSR_384,{COMB_CSR_806,{COMB_CSR_805,{COMB_CSR_804,{COMB_CSR_803,{COMB_CSR_,{COMB_CSR_774,{COMB_CSR_262,{_zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented,_zz_EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented_1}}}}}}}}}} != 32'h00000000);
  assign EU0_CsrAccessPlugin_setup_onDecodeWrite = EU0_CsrAccessPlugin_logic_fsm_startLogic_csrWrite;
  assign EU0_CsrAccessPlugin_setup_onDecodeRead = EU0_CsrAccessPlugin_logic_fsm_startLogic_csrRead;
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_trap = ((! EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented) || EU0_CsrAccessPlugin_setup_onDecodeTrap);
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_write = ((EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL && (! EU0_CsrAccessPlugin_logic_fsm_startLogic_trap)) && EU0_CsrAccessPlugin_logic_fsm_startLogic_csrWrite);
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_read = ((EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL && (! EU0_CsrAccessPlugin_logic_fsm_startLogic_trap)) && EU0_CsrAccessPlugin_logic_fsm_startLogic_csrRead);
  assign EU0_CsrAccessPlugin_setup_onDecodeAddress = _zz_EU0_CsrAccessPlugin_setup_onDecodeAddress[31 : 20];
  assign EU0_CsrAccessPlugin_logic_fsm_startLogic_onDecodeDo = (EU0_ExecutionUnitBase_pipeline_execute_0_valid && EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL);
  assign when_CsrAccessPlugin_l181 = (EU0_CsrAccessPlugin_logic_fsm_startLogic_onDecodeDo && COMB_CSR_384);
  assign EU0_CsrAccessPlugin_setup_onReadAddress = _zz_EU0_CsrAccessPlugin_setup_onReadAddress[31 : 20];
  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = EU0_CsrAccessPlugin_logic_fsm_regs_read;
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        if(when_CsrAccessPlugin_l283) begin
          EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = EU0_CsrAccessPlugin_logic_fsm_regs_read;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign EU0_CsrAccessPlugin_setup_onReadMovingOff = ((! EU0_CsrAccessPlugin_setup_onReadHalt) || EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed);
  assign _zz_322 = zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue(1'b0);
  always @(*) _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue = _zz_322;
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1[31 : 0] = 32'h40141101;
  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2[31 : 31] = PrivilegedPlugin_logic_machine_cause_interrupt;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2[3 : 0] = PrivilegedPlugin_logic_machine_cause_code;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[12 : 11] = PrivilegedPlugin_logic_machine_mstatus_mpp;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[7 : 7] = PrivilegedPlugin_logic_machine_mstatus_mpie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[3 : 3] = PrivilegedPlugin_logic_machine_mstatus_mie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[31 : 31] = PrivilegedPlugin_logic_machine_mstatus_sd;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[14 : 13] = PrivilegedPlugin_logic_machine_mstatus_fs;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[8 : 8] = PrivilegedPlugin_logic_supervisor_sstatus_spp;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[5 : 5] = PrivilegedPlugin_logic_supervisor_sstatus_spie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[1 : 1] = PrivilegedPlugin_logic_supervisor_sstatus_sie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[19 : 19] = MmuPlugin_logic_status_mxr;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[18 : 18] = MmuPlugin_logic_status_sum;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3[17 : 17] = MmuPlugin_logic_status_mprv;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[11 : 11] = PrivilegedPlugin_logic_machine_mip_meip;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[7 : 7] = PrivilegedPlugin_logic_machine_mip_mtip;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[3 : 3] = PrivilegedPlugin_logic_machine_mip_msip;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[9 : 9] = PrivilegedPlugin_logic_supervisor_sip_seipOr;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[5 : 5] = PrivilegedPlugin_logic_supervisor_sip_stip;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4[1 : 1] = PrivilegedPlugin_logic_supervisor_sip_ssip;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[11 : 11] = PrivilegedPlugin_logic_machine_mie_meie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[7 : 7] = PrivilegedPlugin_logic_machine_mie_mtie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[3 : 3] = PrivilegedPlugin_logic_machine_mie_msie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[9 : 9] = PrivilegedPlugin_logic_supervisor_sie_seie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[5 : 5] = PrivilegedPlugin_logic_supervisor_sie_stie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5[1 : 1] = PrivilegedPlugin_logic_supervisor_sie_ssie;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[0 : 0] = PrivilegedPlugin_logic_machine_medeleg_iam;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[3 : 3] = PrivilegedPlugin_logic_machine_medeleg_bp;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[8 : 8] = PrivilegedPlugin_logic_machine_medeleg_eu;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[9 : 9] = PrivilegedPlugin_logic_machine_medeleg_es;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[12 : 12] = PrivilegedPlugin_logic_machine_medeleg_ipf;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[13 : 13] = PrivilegedPlugin_logic_machine_medeleg_lpf;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6[15 : 15] = PrivilegedPlugin_logic_machine_medeleg_spf;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7[9 : 9] = PrivilegedPlugin_logic_machine_mideleg_se;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7[5 : 5] = PrivilegedPlugin_logic_machine_mideleg_st;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7[1 : 1] = PrivilegedPlugin_logic_machine_mideleg_ss;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8[31 : 31] = PrivilegedPlugin_logic_supervisor_cause_interrupt;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8[3 : 0] = PrivilegedPlugin_logic_supervisor_cause_code;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[8 : 8] = PrivilegedPlugin_logic_supervisor_sstatus_spp;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[5 : 5] = PrivilegedPlugin_logic_supervisor_sstatus_spie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[1 : 1] = PrivilegedPlugin_logic_supervisor_sstatus_sie;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[14 : 13] = PrivilegedPlugin_logic_machine_mstatus_fs;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[31 : 31] = PrivilegedPlugin_logic_machine_mstatus_sd;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[19 : 19] = MmuPlugin_logic_status_mxr;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9[18 : 18] = MmuPlugin_logic_status_sum;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10[9 : 9] = (PrivilegedPlugin_logic_supervisor_sie_seie && PrivilegedPlugin_logic_machine_mideleg_se);
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10[5 : 5] = (PrivilegedPlugin_logic_supervisor_sie_stie && PrivilegedPlugin_logic_machine_mideleg_st);
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10[1 : 1] = (PrivilegedPlugin_logic_supervisor_sie_ssie && PrivilegedPlugin_logic_machine_mideleg_ss);
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11[9 : 9] = (PrivilegedPlugin_logic_supervisor_sip_seipOr && PrivilegedPlugin_logic_machine_mideleg_se);
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11[5 : 5] = (PrivilegedPlugin_logic_supervisor_sip_stip && PrivilegedPlugin_logic_machine_mideleg_st);
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11[1 : 1] = (PrivilegedPlugin_logic_supervisor_sip_ssip && PrivilegedPlugin_logic_machine_mideleg_ss);
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12[2 : 0] = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_7;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13[2 : 0] = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_8;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14[2 : 0] = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_9;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15[2 : 0] = _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_10;
  end

  always @(*) begin
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 = 32'h00000000;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16[31 : 31] = MmuPlugin_logic_satp_mode;
    _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16[19 : 0] = MmuPlugin_logic_satp_ppn;
  end

  assign when_CsrAccessPlugin_l244 = (EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_PerformanceCounterPlugin_logic_csrFilter);
  assign _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17[31 : 0] = _zz__zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17;
  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue = (((((_zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 | _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21) | (_zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23 | _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26)) | ((_zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29 | _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31) | (_zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33 | _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35))) | (((_zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37 | _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39) | (_zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41 | _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43)) | ((_zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45 | _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47) | (_zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49 | _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51)))) | ((((REG_CSR_804 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53) | (REG_CSR_805 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54)) | ((REG_CSR_806 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55) | (REG_CSR_384 ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 : _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56))) | (REG_CSR_PerformanceCounterPlugin_logic_csrFilter ? _zz_EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 : 32'h00000000)));
    if(EU0_CsrAccessPlugin_logic_fsm_regs_ramSel) begin
      EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue = EU0_CsrAccessPlugin_logic_ramReadPort_data;
    end
  end

  assign EU0_CsrAccessPlugin_logic_ramReadPort_valid = (EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && EU0_CsrAccessPlugin_logic_fsm_regs_ramSel);
  assign EU0_CsrAccessPlugin_logic_ramReadPort_address = EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress;
  assign when_CsrAccessPlugin_l270 = (EU0_CsrAccessPlugin_logic_ramReadPort_valid && (! EU0_CsrAccessPlugin_logic_ramReadPort_ready));
  always @(*) begin
    EU0_CsrAccessPlugin_setup_onReadToWriteBits = EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
    if(when_CsrAccessPlugin_l276) begin
      EU0_CsrAccessPlugin_setup_onReadToWriteBits[9 : 9] = PrivilegedPlugin_logic_supervisor_sip_seipSoft;
    end
  end

  assign when_CsrAccessPlugin_l276 = (EU0_CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_836);
  assign EU0_CsrAccessPlugin_setup_onWriteMovingOff = ((! EU0_CsrAccessPlugin_setup_onWriteHalt) || EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed);
  assign EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = (EU0_CsrAccessPlugin_logic_fsm_regs_doImm ? _zz_EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask : EU0_CsrAccessPlugin_logic_fsm_regs_rs1);
  assign EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_masked = (EU0_CsrAccessPlugin_logic_fsm_regs_doClear ? (EU0_CsrAccessPlugin_logic_fsm_regs_aluInput & (~ EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask)) : (EU0_CsrAccessPlugin_logic_fsm_regs_aluInput | EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask));
  assign EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_result = (EU0_CsrAccessPlugin_logic_fsm_regs_doMask ? EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_masked : EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask);
  assign EU0_CsrAccessPlugin_setup_onWriteBits = EU0_CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
  assign EU0_CsrAccessPlugin_setup_onWriteAddress = _zz_EU0_CsrAccessPlugin_setup_onWriteAddress[31 : 20];
  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = EU0_CsrAccessPlugin_logic_fsm_regs_write;
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        if(when_CsrAccessPlugin_l309) begin
          EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = EU0_CsrAccessPlugin_logic_fsm_regs_write;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign when_CsrAccessPlugin_l326 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_834);
  assign when_CsrAccessPlugin_l326_1 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_768);
  assign when_CsrAccessPlugin_l326_2 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_836);
  assign when_CsrAccessPlugin_l326_3 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_772);
  assign when_CsrAccessPlugin_l326_4 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_770);
  assign when_CsrAccessPlugin_l326_5 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_771);
  assign when_CsrAccessPlugin_l326_6 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_322);
  assign when_CsrAccessPlugin_l326_7 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_256);
  assign when_CsrAccessPlugin_l326_8 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_260);
  assign when_CsrAccessPlugin_l326_9 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_324);
  assign when_CsrAccessPlugin_l326_10 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_803);
  assign when_CsrAccessPlugin_l326_11 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_804);
  assign when_CsrAccessPlugin_l326_12 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_805);
  assign when_CsrAccessPlugin_l326_13 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_806);
  assign when_CsrAccessPlugin_l331 = ((((MmuPlugin_logic_satpModeWrite != 1'b0) && (MmuPlugin_logic_satpModeWrite != 1'b1)) != 1'b0) == 1'b0);
  assign when_CsrAccessPlugin_l326_14 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_384);
  assign when_CsrAccessPlugin_l325 = (EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PerformanceCounterPlugin_logic_csrFilter);
  assign when_PerformanceCounterPlugin_l273 = (! PerformanceCounterPlugin_logic_csrWrite_fired);
  assign when_PerformanceCounterPlugin_l275 = (! PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready);
  assign when_CsrAccessPlugin_l336 = (EU0_CsrAccessPlugin_logic_ramWritePort_valid && EU0_CsrAccessPlugin_logic_ramWritePort_ready);
  assign EU0_CsrAccessPlugin_logic_ramWritePort_valid = ((EU0_CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && EU0_CsrAccessPlugin_logic_fsm_regs_ramSel) && (! EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired));
  assign EU0_CsrAccessPlugin_logic_ramWritePort_address = EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress;
  assign EU0_CsrAccessPlugin_logic_ramWritePort_data = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign when_CsrAccessPlugin_l340 = (EU0_CsrAccessPlugin_logic_ramWritePort_valid && (! EU0_CsrAccessPlugin_logic_ramWritePort_ready));
  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_isDone = 1'b0;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
        EU0_CsrAccessPlugin_logic_fsm_isDone = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_isCompletionReady = 1'b0;
    if(EU0_ExecutionUnitBase_pipeline_execute_2_ready) begin
      EU0_CsrAccessPlugin_logic_fsm_isCompletionReady = 1'b1;
    end
  end

  always @(*) begin
    EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_stateReg;
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
        if(EU0_CsrAccessPlugin_logic_fsm_startLogic_onDecodeDo) begin
          EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_READ;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        if(when_CsrAccessPlugin_l283) begin
          EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        if(when_CsrAccessPlugin_l309) begin
          EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
        if(EU0_CsrAccessPlugin_logic_fsm_isCompletionReady) begin
          EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed) begin
      EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE;
    end
    if(EU0_CsrAccessPlugin_logic_fsm_wantStart) begin
      EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE;
    end
    if(EU0_CsrAccessPlugin_logic_fsm_wantKill) begin
      EU0_CsrAccessPlugin_logic_fsm_stateNext = EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT;
    end
  end

  assign switch_CsrAccessPlugin_l204 = EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP[31 : 20];
  assign when_CsrAccessPlugin_l283 = (! EU0_CsrAccessPlugin_setup_onReadHalt);
  assign when_CsrAccessPlugin_l309 = (! EU0_CsrAccessPlugin_setup_onWriteHalt);
  assign EU0_CsrAccessPlugin_setup_intFormatPort_payload = EU0_CsrAccessPlugin_logic_fsm_regs_csrValue;
  assign EU0_CsrAccessPlugin_setup_trap_valid = (((EU0_ExecutionUnitBase_pipeline_execute_2_valid && EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL) && EU0_CsrAccessPlugin_logic_fsm_isDone) && (EU0_CsrAccessPlugin_logic_fsm_regs_trap || EU0_CsrAccessPlugin_logic_fsm_regs_flushPipeline));
  assign EU0_CsrAccessPlugin_setup_trap_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  always @(*) begin
    EU0_CsrAccessPlugin_setup_trap_payload_cause = 4'b0010;
    if(when_CsrAccessPlugin_l376) begin
      EU0_CsrAccessPlugin_setup_trap_payload_cause = 4'b1001;
    end
  end

  assign EU0_CsrAccessPlugin_setup_trap_payload_tval = EU0_CsrAccessPlugin_logic_fsm_regs_microOp;
  assign EU0_CsrAccessPlugin_setup_trap_payload_skipCommit = EU0_CsrAccessPlugin_logic_fsm_regs_trap;
  assign EU0_CsrAccessPlugin_setup_trap_payload_reason = 8'h01;
  assign EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_CsrAccessPlugin_l373 = ((EU0_ExecutionUnitBase_pipeline_execute_2_valid && EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL) && (! EU0_CsrAccessPlugin_logic_fsm_isDone));
  assign when_CsrAccessPlugin_l376 = (! EU0_CsrAccessPlugin_logic_fsm_regs_trap);
  assign EU0_ExecutionUnitBase_pipeline_execute_2_isFireing = (EU0_ExecutionUnitBase_pipeline_execute_2_valid && EU0_ExecutionUnitBase_pipeline_execute_2_ready);
  assign csrAccess_valid = ((EU0_ExecutionUnitBase_pipeline_execute_2_isFireing && EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL) && (! EU0_CsrAccessPlugin_logic_fsm_regs_trap));
  assign csrAccess_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  assign csrAccess_payload_address = _zz_csrAccess_payload_address[31 : 20];
  assign csrAccess_payload_write = EU0_CsrAccessPlugin_setup_onWriteBits;
  assign csrAccess_payload_read = EU0_CsrAccessPlugin_logic_fsm_regs_csrValue;
  assign csrAccess_payload_writeDone = EU0_CsrAccessPlugin_logic_fsm_regs_write;
  assign csrAccess_payload_readDone = EU0_CsrAccessPlugin_logic_fsm_regs_read;
  assign DecoderPlugin_logic_slots_0_rdZero = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[11 : 7] == 5'h00);
  assign FrontendPlugin_decoded_LEGAL_0 = ((|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000005f) == 32'h00000017),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000007f) == 32'h0000006f),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & _zz_FrontendPlugin_decoded_LEGAL_0) == 32'h00001073),{(_zz_FrontendPlugin_decoded_LEGAL_0_1 == _zz_FrontendPlugin_decoded_LEGAL_0_2),{_zz_FrontendPlugin_decoded_LEGAL_0_3,{_zz_FrontendPlugin_decoded_LEGAL_0_4,_zz_FrontendPlugin_decoded_LEGAL_0_5}}}}}}) && (! FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_0));
  assign FrontendPlugin_decoded_READ_RS_0_0 = _zz_FrontendPlugin_decoded_READ_RS_0_0[0];
  assign _zz_FrontendPlugin_decoded_SQ_ALLOC_0 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h10000070) == 32'h00000020);
  assign _zz_FrontendPlugin_decoded_SQ_ALLOC_0_1 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h08000070) == 32'h08000020);
  assign FrontendPlugin_decoded_READ_RS_1_0 = _zz_FrontendPlugin_decoded_READ_RS_1_0[0];
  assign _zz_323 = zz_DecoderPlugin_logic_slots_0_x0AlwaysZero(1'b0);
  always @(*) DecoderPlugin_logic_slots_0_x0AlwaysZero = _zz_323;
  assign _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_0 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h0000000c) == 32'h00000004);
  assign _zz_FrontendPlugin_decoded_WRITE_RD_0 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000048) == 32'h00000048);
  assign FrontendPlugin_decoded_WRITE_RD_0 = (_zz_FrontendPlugin_decoded_WRITE_RD_0_1[0] && (! (DecoderPlugin_logic_slots_0_rdZero && DecoderPlugin_logic_slots_0_x0AlwaysZero)));
  assign _zz_FrontendPlugin_decoded_IS_ANY_0 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 & 32'h00000050) == 32'h00000040);
  assign FrontendPlugin_decoded_ALU0_ALU1_SEL_0 = _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_0_1[0];
  assign FrontendPlugin_decoded_EU0_SEL_0 = _zz_FrontendPlugin_decoded_EU0_SEL_0[0];
  assign FrontendPlugin_decoded_LQ_ALLOC_0 = _zz_FrontendPlugin_decoded_LQ_ALLOC_0[0];
  assign FrontendPlugin_decoded_SQ_ALLOC_0 = _zz_FrontendPlugin_decoded_SQ_ALLOC_0_2[0];
  assign FrontendPlugin_decoded_TRAP_0 = (FrontendPlugin_decoded_Frontend_MASK_ALIGNED_0 && ((((! FrontendPlugin_decoded_LEGAL_0) || FrontendPlugin_decoded_Frontend_FETCH_FAULT_0) || DecoderPlugin_setup_trapRaise) || DecoderPlugin_setup_debugEnter_0));
  assign FrontendPlugin_decoded_Frontend_DECODED_MASK_0 = (FrontendPlugin_decoded_Frontend_MASK_ALIGNED_0 && (! (FrontendPlugin_decoded_TRAP_0 != 1'b0)));
  assign FrontendPlugin_decoded_Frontend_MICRO_OP_0 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0;
  assign FrontendPlugin_decoded_ARCH_RD_0 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[11 : 7];
  assign FrontendPlugin_decoded_ARCH_RS_0_0 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[19 : 15];
  assign FrontendPlugin_decoded_ARCH_RS_1_0 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[24 : 20];
  assign DecoderPlugin_logic_slots_1_rdZero = (FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[11 : 7] == 5'h00);
  assign FrontendPlugin_decoded_LEGAL_1 = ((|{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000005f) == 32'h00000017),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000007f) == 32'h0000006f),{((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & _zz_FrontendPlugin_decoded_LEGAL_1) == 32'h00001073),{(_zz_FrontendPlugin_decoded_LEGAL_1_1 == _zz_FrontendPlugin_decoded_LEGAL_1_2),{_zz_FrontendPlugin_decoded_LEGAL_1_3,{_zz_FrontendPlugin_decoded_LEGAL_1_4,_zz_FrontendPlugin_decoded_LEGAL_1_5}}}}}}) && (! FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_1));
  assign FrontendPlugin_decoded_READ_RS_0_1 = _zz_FrontendPlugin_decoded_READ_RS_0_1[0];
  assign _zz_FrontendPlugin_decoded_SQ_ALLOC_1 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h10000070) == 32'h00000020);
  assign _zz_FrontendPlugin_decoded_SQ_ALLOC_1_1 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h08000070) == 32'h08000020);
  assign FrontendPlugin_decoded_READ_RS_1_1 = _zz_FrontendPlugin_decoded_READ_RS_1_1[0];
  assign _zz_324 = zz_DecoderPlugin_logic_slots_1_x0AlwaysZero(1'b0);
  always @(*) DecoderPlugin_logic_slots_1_x0AlwaysZero = _zz_324;
  assign _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_1 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h0000000c) == 32'h00000004);
  assign _zz_FrontendPlugin_decoded_IS_JAL_1 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000048) == 32'h00000048);
  assign FrontendPlugin_decoded_WRITE_RD_1 = (_zz_FrontendPlugin_decoded_WRITE_RD_1[0] && (! (DecoderPlugin_logic_slots_1_rdZero && DecoderPlugin_logic_slots_1_x0AlwaysZero)));
  assign _zz_FrontendPlugin_decoded_IS_ANY_1 = ((FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 & 32'h00000050) == 32'h00000040);
  assign FrontendPlugin_decoded_ALU0_ALU1_SEL_1 = _zz_FrontendPlugin_decoded_ALU0_ALU1_SEL_1_1[0];
  assign FrontendPlugin_decoded_EU0_SEL_1 = _zz_FrontendPlugin_decoded_EU0_SEL_1[0];
  assign FrontendPlugin_decoded_LQ_ALLOC_1 = _zz_FrontendPlugin_decoded_LQ_ALLOC_1[0];
  assign FrontendPlugin_decoded_SQ_ALLOC_1 = _zz_FrontendPlugin_decoded_SQ_ALLOC_1_2[0];
  assign FrontendPlugin_decoded_TRAP_1 = (FrontendPlugin_decoded_Frontend_MASK_ALIGNED_1 && ((((! FrontendPlugin_decoded_LEGAL_1) || FrontendPlugin_decoded_Frontend_FETCH_FAULT_1) || DecoderPlugin_setup_trapRaise) || DecoderPlugin_setup_debugEnter_1));
  assign FrontendPlugin_decoded_Frontend_DECODED_MASK_1 = (FrontendPlugin_decoded_Frontend_MASK_ALIGNED_1 && (! ({FrontendPlugin_decoded_TRAP_1,FrontendPlugin_decoded_TRAP_0} != 2'b00)));
  assign FrontendPlugin_decoded_Frontend_MICRO_OP_1 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1;
  assign FrontendPlugin_decoded_ARCH_RD_1 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[11 : 7];
  assign FrontendPlugin_decoded_ARCH_RS_0_1 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[19 : 15];
  assign FrontendPlugin_decoded_ARCH_RS_1_1 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[24 : 20];
  assign DecoderPlugin_logic_exception_set = (FrontendPlugin_decoded_isFireing && ({FrontendPlugin_decoded_TRAP_1,FrontendPlugin_decoded_TRAP_0} != 2'b00));
  assign DecoderPlugin_logic_exception_clear = FrontendPlugin_decoded_isFlushed;
  assign when_DecoderPlugin_l302 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l303 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l304 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l306 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l307 = (! DecoderPlugin_logic_exception_trigged);
  assign when_DecoderPlugin_l308 = (! DecoderPlugin_logic_exception_trigged);
  assign _zz_DecoderPlugin_setup_exceptionPort_payload_tval = {DecoderPlugin_logic_exception_exceptionReg_1,DecoderPlugin_logic_exception_exceptionReg_0};
  assign _zz_DecoderPlugin_setup_exceptionPort_payload_tval_1 = _zz__zz_DecoderPlugin_setup_exceptionPort_payload_tval_1[1];
  assign DecoderPlugin_logic_exception_fetchFault = _zz_DecoderPlugin_logic_exception_fetchFault[0];
  assign DecoderPlugin_logic_exception_fetchFaultPage = _zz_DecoderPlugin_logic_exception_fetchFaultPage[0];
  assign DecoderPlugin_logic_exception_debugEnter = _zz_DecoderPlugin_logic_exception_debugEnter[0];
  assign DecoderPlugin_logic_exception_pc = ((DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_epcReg_0 : 32'h00000000) | (_zz_DecoderPlugin_setup_exceptionPort_payload_tval_1 ? DecoderPlugin_logic_exception_epcReg_1 : 32'h00000000));
  assign DecoderPlugin_logic_exception_pipelineEmpty = ((! FrontendPlugin_isBusyAfterDecode) && CommitPlugin_setup_isRobEmpty);
  assign DecoderPlugin_logic_exception_doIt = (DecoderPlugin_logic_exception_trigged && DecoderPlugin_logic_exception_pipelineEmpty);
  assign _zz_FrontendPlugin_decoded_isFlushingRoot = (DecoderPlugin_logic_exception_doIt || DecoderPlugin_logic_exception_doItAgain);
  assign FrontendPlugin_decoded_haltRequest_DecoderPlugin_l322 = DecoderPlugin_logic_exception_trigged;
  assign FrontendPlugin_decoded_haltRequest_DecoderPlugin_l323 = (DecoderPlugin_setup_trapHalt && (! DecoderPlugin_setup_trapRaise));
  assign DecoderPlugin_setup_trapReady = (FrontendPlugin_decoded_valid && DecoderPlugin_logic_exception_pipelineEmpty);
  assign DecoderPlugin_setup_exceptionPort_valid = DecoderPlugin_logic_exception_doIt;
  assign DecoderPlugin_setup_exceptionPort_payload_epc = DecoderPlugin_logic_exception_pc;
  always @(*) begin
    if(DecoderPlugin_logic_exception_fetchFault) begin
      if(DecoderPlugin_logic_exception_fetchFaultPage) begin
        DecoderPlugin_setup_exceptionPort_payload_cause = 4'b1100;
      end else begin
        DecoderPlugin_setup_exceptionPort_payload_cause = 4'b0001;
      end
    end else begin
      DecoderPlugin_setup_exceptionPort_payload_cause = 4'b0010;
    end
  end

  always @(*) begin
    if(DecoderPlugin_logic_exception_fetchFault) begin
      DecoderPlugin_setup_exceptionPort_payload_tval = _zz_DecoderPlugin_setup_exceptionPort_payload_tval_2;
    end else begin
      DecoderPlugin_setup_exceptionPort_payload_tval = ((DecoderPlugin_logic_exception_exceptionReg_0 ? DecoderPlugin_logic_exception_instReg_0 : 32'h00000000) | (_zz_DecoderPlugin_setup_exceptionPort_payload_tval_1 ? DecoderPlugin_logic_exception_instReg_1 : 32'h00000000));
    end
  end

  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h00001048) == 32'h00001008);
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h00002050) == 32'h00002050);
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_1 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h02000050) == 32'h02000050);
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_1 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_0 & 32'h00001050) == 32'h00001050);
  assign FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0_2[0];
  assign FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0_2[0];
  assign FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0 = _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_0[0];
  assign FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0[0];
  assign FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0[0];
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_1 & 32'h00001048) == 32'h00001008);
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_1 & 32'h00002050) == 32'h00002050);
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_1 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_1 & 32'h02000050) == 32'h02000050);
  assign _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_1 = ((FrontendPlugin_serialized_Frontend_MICRO_OP_1 & 32'h00001050) == 32'h00001050);
  assign FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1_2[0];
  assign FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1 = _zz_FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1_2[0];
  assign FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_1 = _zz_FrontendPlugin_serialized_DispatchPlugin_SPARSE_ROB_LINE_1[0];
  assign FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_1 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_1[0];
  assign FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_1 = _zz_FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_1[0];
  assign FrontendPlugin_dispatch_LATENCY_0_0 = (|{((FrontendPlugin_dispatch_Frontend_MICRO_OP_0 & 32'h00000048) == 32'h00000048),{((FrontendPlugin_dispatch_Frontend_MICRO_OP_0 & 32'h00000030) == 32'h00000010),{((FrontendPlugin_dispatch_Frontend_MICRO_OP_0 & 32'h0000000c) == 32'h00000004),((FrontendPlugin_dispatch_Frontend_MICRO_OP_0 & 32'h02000050) == 32'h00000010)}}});
  assign FrontendPlugin_dispatch_LATENCY_0_1 = (|{((FrontendPlugin_dispatch_Frontend_MICRO_OP_1 & 32'h00000048) == 32'h00000048),{((FrontendPlugin_dispatch_Frontend_MICRO_OP_1 & 32'h00000030) == 32'h00000010),{((FrontendPlugin_dispatch_Frontend_MICRO_OP_1 & 32'h0000000c) == 32'h00000004),((FrontendPlugin_dispatch_Frontend_MICRO_OP_1 & 32'h02000050) == 32'h00000010)}}});
  assign FrontendPlugin_decoded_IS_JAL_0 = _zz_FrontendPlugin_decoded_IS_JAL_0[0];
  assign FrontendPlugin_decoded_IS_JALR_0 = _zz_FrontendPlugin_decoded_IS_JALR_0[0];
  assign FrontendPlugin_decoded_Prediction_IS_BRANCH_0 = _zz_FrontendPlugin_decoded_Prediction_IS_BRANCH_0[0];
  assign FrontendPlugin_decoded_IS_ANY_0 = _zz_FrontendPlugin_decoded_IS_ANY_0_1[0];
  assign switch_Misc_l232_3 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0[2];
  always @(*) begin
    case(switch_Misc_l232_3)
      1'b0 : begin
        _zz_FrontendPlugin_decoded_OFFSET_0 = {{19{_zz__zz_FrontendPlugin_decoded_OFFSET_0[12]}}, _zz__zz_FrontendPlugin_decoded_OFFSET_0};
      end
      default : begin
        _zz_FrontendPlugin_decoded_OFFSET_0 = {{11{_zz__zz_FrontendPlugin_decoded_OFFSET_0_1[20]}}, _zz__zz_FrontendPlugin_decoded_OFFSET_0_1};
      end
    endcase
  end

  assign FrontendPlugin_decoded_OFFSET_0 = _zz_FrontendPlugin_decoded_OFFSET_0;
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink = ({(FrontendPlugin_decoded_ARCH_RD_0 == 5'h05),(FrontendPlugin_decoded_ARCH_RD_0 == 5'h01)} != 2'b00);
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rs1Link = ({(FrontendPlugin_decoded_ARCH_RS_0_0 == 5'h05),(FrontendPlugin_decoded_ARCH_RS_0_0 == 5'h01)} != 2'b00);
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdEquRs1 = (FrontendPlugin_decoded_ARCH_RD_0 == FrontendPlugin_decoded_ARCH_RS_0_0);
  assign FrontendPlugin_decoded_RAS_PUSH_0 = ((FrontendPlugin_decoded_IS_JAL_0 || FrontendPlugin_decoded_IS_JALR_0) && DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink);
  assign FrontendPlugin_decoded_RAS_POP_0 = (FrontendPlugin_decoded_IS_JALR_0 && (((! DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink) && DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rs1Link) || ((DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdLink && DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rs1Link) && (! DecoderPredictionPlugin_logic_decodePatch_slots_0_decode_rdEquRs1))));
  assign FrontendPlugin_decoded_LAST_SLICE_0 = (FrontendPlugin_decoded_PC_0[2 : 2] + 1'b0);
  assign FrontendPlugin_decoded_CONDITIONAL_PREDICTION_0 = FrontendPlugin_decoded_Prediction_CONDITIONAL_TAKE_IT_0[FrontendPlugin_decoded_LAST_SLICE_0];
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices = (_zz_DecoderPredictionPlugin_logic_decodePatch_slots_0_pcAdd_slices + {1'b0,1'b1});
  assign FrontendPlugin_decoded_PC_INC_0 = _zz_FrontendPlugin_decoded_PC_INC_0;
  assign FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0 = ($signed(_zz_FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0) + $signed(FrontendPlugin_decoded_OFFSET_0));
  assign FrontendPlugin_decoded_BAD_RET_PC_0 = (FrontendPlugin_decoded_RAS_POP_0 && (DecoderPredictionPlugin_logic_ras_read != FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_0));
  assign FrontendPlugin_decoded_CAN_IMPROVE_0 = ((! FrontendPlugin_decoded_IS_JALR_0) || FrontendPlugin_decoded_RAS_POP_0);
  assign FrontendPlugin_decoded_BRANCHED_PREDICTION_0 = (((FrontendPlugin_decoded_Prediction_IS_BRANCH_0 && FrontendPlugin_decoded_CONDITIONAL_PREDICTION_0) || FrontendPlugin_decoded_IS_JAL_0) || FrontendPlugin_decoded_IS_JALR_0);
  always @(*) begin
    FrontendPlugin_serialized_PC_TARGET_0 = FrontendPlugin_serialized_PC_TARGET_PRE_RAS_0;
    if(FrontendPlugin_serialized_IS_JALR_0) begin
      FrontendPlugin_serialized_PC_TARGET_0 = DecoderPredictionPlugin_logic_ras_read;
    end
  end

  assign FrontendPlugin_serialized_PC_PREDICTION_0 = (FrontendPlugin_serialized_BRANCHED_PREDICTION_0 ? FrontendPlugin_serialized_PC_TARGET_0 : FrontendPlugin_serialized_PC_INC_0);
  assign DecoderPredictionPlugin_logic_decodePatch_slots_0_applyIt_badTaken = (FrontendPlugin_serialized_IS_ANY_0 ? (FrontendPlugin_serialized_BRANCHED_PREDICTION_0 != FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0) : FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0);
  assign FrontendPlugin_serialized_MISSMATCH_PC_0 = (DecoderPredictionPlugin_logic_decodePatch_slots_0_applyIt_badTaken || FrontendPlugin_serialized_BAD_RET_PC_0);
  assign FrontendPlugin_serialized_MISSMATCH_HISTORY_0 = 1'b0;
  assign FrontendPlugin_serialized_MISSMATCH_0 = (FrontendPlugin_serialized_MISSMATCH_PC_0 || FrontendPlugin_serialized_MISSMATCH_HISTORY_0);
  assign FrontendPlugin_serialized_NEED_CORRECTION_0 = ((FrontendPlugin_serialized_Frontend_DECODED_MASK_0 && FrontendPlugin_serialized_CAN_IMPROVE_0) && FrontendPlugin_serialized_MISSMATCH_0);
  assign FrontendPlugin_serialized_BRANCH_SEL_0 = FrontendPlugin_serialized_IS_ANY_0;
  always @(*) begin
    if(FrontendPlugin_serialized_NEED_CORRECTION_0) begin
      FrontendPlugin_serialized_BRANCH_EARLY_0_taken = FrontendPlugin_serialized_BRANCHED_PREDICTION_0;
    end else begin
      FrontendPlugin_serialized_BRANCH_EARLY_0_taken = FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0;
    end
  end

  always @(*) begin
    if(FrontendPlugin_serialized_NEED_CORRECTION_0) begin
      FrontendPlugin_serialized_BRANCH_EARLY_0_pc = FrontendPlugin_serialized_PC_TARGET_0;
    end else begin
      FrontendPlugin_serialized_BRANCH_EARLY_0_pc = FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
    end
  end

  assign when_DecoderPredictionPlugin_l212 = (FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0 && FrontendPlugin_serialized_RAS_PUSH_0);
  assign when_DecoderPredictionPlugin_l213 = (! DecoderPredictionPlugin_logic_decodePatch_rasPushUsed);
  assign when_DecoderPredictionPlugin_l219 = (FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0 && FrontendPlugin_serialized_RAS_POP_0);
  assign FrontendPlugin_serialized_DecoderPredictionPlugin_RAS_PUSH_PTR_0 = DecoderPredictionPlugin_logic_ras_ptr_push;
  assign FrontendPlugin_decoded_IS_JAL_1 = _zz_FrontendPlugin_decoded_IS_JAL_1_1[0];
  assign FrontendPlugin_decoded_IS_JALR_1 = _zz_FrontendPlugin_decoded_IS_JALR_1[0];
  assign FrontendPlugin_decoded_Prediction_IS_BRANCH_1 = _zz_FrontendPlugin_decoded_Prediction_IS_BRANCH_1[0];
  assign FrontendPlugin_decoded_IS_ANY_1 = _zz_FrontendPlugin_decoded_IS_ANY_1_1[0];
  assign switch_Misc_l232_4 = FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1[2];
  always @(*) begin
    case(switch_Misc_l232_4)
      1'b0 : begin
        _zz_FrontendPlugin_decoded_OFFSET_1 = {{19{_zz__zz_FrontendPlugin_decoded_OFFSET_1[12]}}, _zz__zz_FrontendPlugin_decoded_OFFSET_1};
      end
      default : begin
        _zz_FrontendPlugin_decoded_OFFSET_1 = {{11{_zz__zz_FrontendPlugin_decoded_OFFSET_1_1[20]}}, _zz__zz_FrontendPlugin_decoded_OFFSET_1_1};
      end
    endcase
  end

  assign FrontendPlugin_decoded_OFFSET_1 = _zz_FrontendPlugin_decoded_OFFSET_1;
  assign DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rdLink = ({(FrontendPlugin_decoded_ARCH_RD_1 == 5'h05),(FrontendPlugin_decoded_ARCH_RD_1 == 5'h01)} != 2'b00);
  assign DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rs1Link = ({(FrontendPlugin_decoded_ARCH_RS_0_1 == 5'h05),(FrontendPlugin_decoded_ARCH_RS_0_1 == 5'h01)} != 2'b00);
  assign DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rdEquRs1 = (FrontendPlugin_decoded_ARCH_RD_1 == FrontendPlugin_decoded_ARCH_RS_0_1);
  assign FrontendPlugin_decoded_RAS_PUSH_1 = ((FrontendPlugin_decoded_IS_JAL_1 || FrontendPlugin_decoded_IS_JALR_1) && DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rdLink);
  assign FrontendPlugin_decoded_RAS_POP_1 = (FrontendPlugin_decoded_IS_JALR_1 && (((! DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rdLink) && DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rs1Link) || ((DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rdLink && DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rs1Link) && (! DecoderPredictionPlugin_logic_decodePatch_slots_1_decode_rdEquRs1))));
  assign FrontendPlugin_decoded_LAST_SLICE_1 = (FrontendPlugin_decoded_PC_1[2 : 2] + 1'b0);
  assign FrontendPlugin_decoded_CONDITIONAL_PREDICTION_1 = FrontendPlugin_decoded_Prediction_CONDITIONAL_TAKE_IT_1[FrontendPlugin_decoded_LAST_SLICE_1];
  assign DecoderPredictionPlugin_logic_decodePatch_slots_1_pcAdd_slices = (_zz_DecoderPredictionPlugin_logic_decodePatch_slots_1_pcAdd_slices + {1'b0,1'b1});
  assign FrontendPlugin_decoded_PC_INC_1 = _zz_FrontendPlugin_decoded_PC_INC_1;
  assign FrontendPlugin_decoded_PC_TARGET_PRE_RAS_1 = ($signed(_zz_FrontendPlugin_decoded_PC_TARGET_PRE_RAS_1) + $signed(FrontendPlugin_decoded_OFFSET_1));
  assign FrontendPlugin_decoded_BAD_RET_PC_1 = (FrontendPlugin_decoded_RAS_POP_1 && (DecoderPredictionPlugin_logic_ras_read != FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_1));
  assign FrontendPlugin_decoded_CAN_IMPROVE_1 = ((! FrontendPlugin_decoded_IS_JALR_1) || FrontendPlugin_decoded_RAS_POP_1);
  assign FrontendPlugin_decoded_BRANCHED_PREDICTION_1 = (((FrontendPlugin_decoded_Prediction_IS_BRANCH_1 && FrontendPlugin_decoded_CONDITIONAL_PREDICTION_1) || FrontendPlugin_decoded_IS_JAL_1) || FrontendPlugin_decoded_IS_JALR_1);
  always @(*) begin
    FrontendPlugin_serialized_PC_TARGET_1 = FrontendPlugin_serialized_PC_TARGET_PRE_RAS_1;
    if(FrontendPlugin_serialized_IS_JALR_1) begin
      FrontendPlugin_serialized_PC_TARGET_1 = DecoderPredictionPlugin_logic_ras_read;
    end
  end

  assign FrontendPlugin_serialized_PC_PREDICTION_1 = (FrontendPlugin_serialized_BRANCHED_PREDICTION_1 ? FrontendPlugin_serialized_PC_TARGET_1 : FrontendPlugin_serialized_PC_INC_1);
  assign DecoderPredictionPlugin_logic_decodePatch_slots_1_applyIt_badTaken = (FrontendPlugin_serialized_IS_ANY_1 ? (FrontendPlugin_serialized_BRANCHED_PREDICTION_1 != FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_1) : FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_1);
  assign FrontendPlugin_serialized_MISSMATCH_PC_1 = (DecoderPredictionPlugin_logic_decodePatch_slots_1_applyIt_badTaken || FrontendPlugin_serialized_BAD_RET_PC_1);
  assign FrontendPlugin_serialized_MISSMATCH_HISTORY_1 = 1'b0;
  assign FrontendPlugin_serialized_MISSMATCH_1 = (FrontendPlugin_serialized_MISSMATCH_PC_1 || FrontendPlugin_serialized_MISSMATCH_HISTORY_1);
  assign FrontendPlugin_serialized_NEED_CORRECTION_1 = ((FrontendPlugin_serialized_Frontend_DECODED_MASK_1 && FrontendPlugin_serialized_CAN_IMPROVE_1) && FrontendPlugin_serialized_MISSMATCH_1);
  assign FrontendPlugin_serialized_BRANCH_SEL_1 = FrontendPlugin_serialized_IS_ANY_1;
  always @(*) begin
    if(FrontendPlugin_serialized_NEED_CORRECTION_1) begin
      FrontendPlugin_serialized_BRANCH_EARLY_1_taken = FrontendPlugin_serialized_BRANCHED_PREDICTION_1;
    end else begin
      FrontendPlugin_serialized_BRANCH_EARLY_1_taken = FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_1;
    end
  end

  always @(*) begin
    if(FrontendPlugin_serialized_NEED_CORRECTION_1) begin
      FrontendPlugin_serialized_BRANCH_EARLY_1_pc = FrontendPlugin_serialized_PC_TARGET_1;
    end else begin
      FrontendPlugin_serialized_BRANCH_EARLY_1_pc = FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_PC_NEXT_1;
    end
  end

  assign when_DecoderPredictionPlugin_l212_1 = (FrontendPlugin_serialized_Frontend_DISPATCH_MASK_1 && FrontendPlugin_serialized_RAS_PUSH_1);
  assign when_DecoderPredictionPlugin_l213_1 = (! DecoderPredictionPlugin_logic_decodePatch_rasPushUsed_1);
  assign when_DecoderPredictionPlugin_l219_1 = (FrontendPlugin_serialized_Frontend_DISPATCH_MASK_1 && FrontendPlugin_serialized_RAS_POP_1);
  assign FrontendPlugin_serialized_DecoderPredictionPlugin_RAS_PUSH_PTR_1 = DecoderPredictionPlugin_logic_ras_ptr_push;
  assign DecoderPredictionPlugin_logic_decodePatch_applyIt_hit = ({FrontendPlugin_serialized_NEED_CORRECTION_1,FrontendPlugin_serialized_NEED_CORRECTION_0} != 2'b00);
  assign FrontendPlugin_serialized_isFireing = (FrontendPlugin_serialized_valid && FrontendPlugin_serialized_ready);
  assign when_DecoderPredictionPlugin_l236 = (FrontendPlugin_serialized_ready || FrontendPlugin_serialized_isFlushed);
  assign DecoderPredictionPlugin_setup_decodeJump_valid = (FrontendPlugin_serialized_valid && DecoderPredictionPlugin_logic_decodePatch_applyIt_hit);
  assign DecoderPredictionPlugin_setup_decodeJump_payload_pc = _zz_DecoderPredictionPlugin_setup_decodeJump_payload_pc;
  assign DecoderPredictionPlugin_setup_historyPush_flush = DecoderPredictionPlugin_setup_decodeJump_valid;
  assign when_DecoderPredictionPlugin_l243 = (! FrontendPlugin_serialized_isFireing);
  assign when_DecoderPredictionPlugin_l244 = (! FrontendPlugin_serialized_isFireing);
  assign FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0 = (FrontendPlugin_serialized_Frontend_DECODED_MASK_0 && (! 1'b0));
  assign FrontendPlugin_serialized_Frontend_DISPATCH_MASK_1 = (FrontendPlugin_serialized_Frontend_DECODED_MASK_1 && (! (FrontendPlugin_serialized_NEED_CORRECTION_0 != 1'b0)));
  always @(*) begin
    DecoderPredictionPlugin_setup_historyPush_mask[0] = ((((FrontendPlugin_serialized_valid && DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle) && FrontendPlugin_serialized_Prediction_IS_BRANCH_0) && FrontendPlugin_serialized_Frontend_DECODED_MASK_0) && (! 1'b0));
    DecoderPredictionPlugin_setup_historyPush_mask[1] = ((((FrontendPlugin_serialized_valid && DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle) && FrontendPlugin_serialized_Prediction_IS_BRANCH_1) && FrontendPlugin_serialized_Frontend_DECODED_MASK_1) && (! (FrontendPlugin_serialized_NEED_CORRECTION_0 != 1'b0)));
  end

  always @(*) begin
    DecoderPredictionPlugin_setup_historyPush_taken[0] = FrontendPlugin_serialized_BRANCHED_PREDICTION_0;
    DecoderPredictionPlugin_setup_historyPush_taken[1] = FrontendPlugin_serialized_BRANCHED_PREDICTION_1;
  end

  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_valid = ALU0_ExecutionUnitBase_pipeline_push_port_valid;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID = ALU0_ExecutionUnitBase_pipeline_push_port_robId;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD = ALU0_ExecutionUnitBase_pipeline_push_port_physRd;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1[31 : 0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_1[5 : 0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_1[5 : 0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_PC = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC_1[31 : 0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_1[3 : 0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL = ((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000044) == 32'h00000004);
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1 = {(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004004) == 32'h00004000)),(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00006004) == 32'h00002000))};
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1 = {(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001000) == 32'h00001000)),(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00003000) == 32'h00002000))};
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = ((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000010) == 32'h00000000);
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1[0];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1 = {(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h0000000c) == 32'h00000004)),(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000008) == 32'h00000008))};
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1;
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2 = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO[0];
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC1_CTRL = (|_zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL);
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL = {(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000004) == 32'h00000004)),(|((ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000024) == 32'h00000000))};
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED = _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED[0];
  assign ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid = ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  assign ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address = ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1 = ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  assign ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid = ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  assign ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address = ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2 = ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  assign ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid = ((ALU0_ExecutionUnitBase_pipeline_execute_0_valid && ALU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD) && (ALU0_IntFormatPlugin_logic_stages_0_wb_valid != 1'b0));
  assign ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId = ALU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  assign ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_address = ALU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  assign ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_data = ALU0_IntFormatPlugin_logic_stages_0_wb_payload;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_isFireing = (ALU0_ExecutionUnitBase_pipeline_execute_0_valid && ALU0_ExecutionUnitBase_pipeline_execute_0_ready);
  assign ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid = (ALU0_ExecutionUnitBase_pipeline_execute_0_isFireing && ALU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E0);
  assign ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id = ALU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  assign ALU0_ExecutionUnitBase_pipeline_completion_1_port_valid = (ALU0_ExecutionUnitBase_pipeline_execute_1_isFireing && ALU0_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E1);
  assign ALU0_ExecutionUnitBase_pipeline_completion_1_port_payload_id = ALU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
  assign ALU0_ExecutionUnitBase_pipeline_execute_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU0_ExecutionUnitBase_pipeline_fetch_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ready = 1'b1;
  assign ALU0_ExecutionUnitBase_pipeline_execute_1_ready = 1'b1;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_valid = ALU0_ExecutionUnitBase_pipeline_fetch_1_valid;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2 = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED = ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_SEL = ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_SEL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL = ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL = ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SEL = ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SEL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT = ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_LEFT;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SIGNED = ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SIGNED;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL = ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_SEL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL = ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP = ALU0_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_PC = ALU0_ExecutionUnitBase_pipeline_fetch_1_PC;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID = ALU0_ExecutionUnitBase_pipeline_fetch_1_BRANCH_ID;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD = ALU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID = ALU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD = ALU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E0 = ALU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E0;
  assign ALU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E1 = ALU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E1;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_valid = ALU1_ExecutionUnitBase_pipeline_push_port_valid;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID = ALU1_ExecutionUnitBase_pipeline_push_port_robId;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD = ALU1_ExecutionUnitBase_pipeline_push_port_physRd;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1[31 : 0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0_1[5 : 0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1[0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1_1[5 : 0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1[0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1[0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_PC = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PC_1[31 : 0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID_1[3 : 0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL = ((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000044) == 32'h00000004);
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL_1[0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1 = {(|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00004004) == 32'h00004000)),(|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00006004) == 32'h00002000))};
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_1;
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL_2;
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1 = {(|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001000) == 32'h00001000)),(|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00003000) == 32'h00002000))};
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_1;
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL_2;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL[0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT[0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = ((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000010) == 32'h00000000);
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL[0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1[0];
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1 = {(|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h0000000c) == 32'h00000004)),(|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000008) == 32'h00000008))};
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_1;
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2 = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL_2;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT_1[0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO[0];
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC1_CTRL = (|_zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL);
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL = {(|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000004) == 32'h00000004)),(|((ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000024) == 32'h00000000))};
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED = _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED[0];
  assign ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid = ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  assign ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address = ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_integer_RS1 = ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  assign ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid = ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  assign ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address = ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_integer_RS2 = ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  assign ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_valid = ((ALU1_ExecutionUnitBase_pipeline_execute_0_valid && ALU1_ExecutionUnitBase_pipeline_execute_0_WRITE_RD) && (ALU1_IntFormatPlugin_logic_stages_0_wb_valid != 1'b0));
  assign ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_robId = ALU1_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  assign ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_address = ALU1_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
  assign ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_data = ALU1_IntFormatPlugin_logic_stages_0_wb_payload;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_isFireing = (ALU1_ExecutionUnitBase_pipeline_execute_0_valid && ALU1_ExecutionUnitBase_pipeline_execute_0_ready);
  assign ALU1_ExecutionUnitBase_pipeline_completion_0_port_valid = (ALU1_ExecutionUnitBase_pipeline_execute_0_isFireing && ALU1_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E0);
  assign ALU1_ExecutionUnitBase_pipeline_completion_0_port_payload_id = ALU1_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
  assign ALU1_ExecutionUnitBase_pipeline_completion_1_port_valid = (ALU1_ExecutionUnitBase_pipeline_execute_1_isFireing && ALU1_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E1);
  assign ALU1_ExecutionUnitBase_pipeline_completion_1_port_payload_id = ALU1_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
  assign ALU1_ExecutionUnitBase_pipeline_execute_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU1_ExecutionUnitBase_pipeline_fetch_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_ready = 1'b1;
  assign ALU1_ExecutionUnitBase_pipeline_execute_1_ready = 1'b1;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_valid = ALU1_ExecutionUnitBase_pipeline_fetch_1_valid;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2 = ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT = ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO = ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 = ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_SrcStageables_UNSIGNED = ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_SEL = ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_SEL;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_BITWISE_CTRL = ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_IntAluPlugin_ALU_CTRL = ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SEL = ALU1_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SEL;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_LEFT = ALU1_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_LEFT;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_ShiftPlugin_SIGNED = ALU1_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SIGNED;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL = ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_SEL;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL = ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP = ALU1_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_PC = ALU1_ExecutionUnitBase_pipeline_fetch_1_PC;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID = ALU1_ExecutionUnitBase_pipeline_fetch_1_BRANCH_ID;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_WRITE_RD = ALU1_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_ROB_ID = ALU1_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_PHYS_RD = ALU1_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E0 = ALU1_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E0;
  assign ALU1_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E1 = ALU1_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E1;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_valid = EU0_ExecutionUnitBase_pipeline_push_port_valid;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID = EU0_ExecutionUnitBase_pipeline_push_port_robId;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD = EU0_ExecutionUnitBase_pipeline_push_port_physRd;
  assign EU0_ExecutionUnitBase_pipeline_push_port_ready = EU0_ExecutionUnitBase_pipeline_fetch_0_ready;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0 = EU0_ExecutionUnitBase_pipeline_push_port_context_0;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1 = EU0_ExecutionUnitBase_pipeline_push_port_context_1;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_2[31 : 0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_2[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_2[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_2[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_PC = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_2[31 : 0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_2[4 : 0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_2[0 : 0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2 = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00002000) == 32'h00002000);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00001000) == 32'h00001000);
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00006000) == 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC[0];
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD = ((EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP & 32'h00000020) == 32'h00000000);
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_FLOAT[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_WFI[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR_1[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO = _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO[0];
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_SrcPlugin_logic_SRC2_CTRL = (|_zz_EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD);
  assign EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_valid = EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0;
  assign EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address = EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1 = EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data;
  assign EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_valid = EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1;
  assign EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address = EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2 = EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data;
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid = ((EU0_ExecutionUnitBase_pipeline_execute_2_valid && EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD) && (EU0_IntFormatPlugin_logic_stages_0_wb_valid != 1'b0));
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_address = EU0_ExecutionUnitBase_pipeline_execute_2_PHYS_RD;
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_data = EU0_IntFormatPlugin_logic_stages_0_wb_payload;
  assign EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_ExecutionUnitBase_l303 = (EU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid && (! EU0_ExecutionUnitBase_pipeline_writeBack_0_write_ready));
  assign EU0_ExecutionUnitBase_pipeline_completion_0_port_valid = (EU0_ExecutionUnitBase_pipeline_execute_2_isFireing && EU0_ExecutionUnitBase_pipeline_execute_2_completion_SEL_E2);
  assign EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_fire = (EU0_ExecutionUnitBase_pipeline_execute_2_isFireing && ({EU0_CsrAccessPlugin_logic_wake_wakeRobsSel,{EU0_DivPlugin_logic_wake_wakeRobsSel,EU0_MulPlugin_logic_wake_wakeRobsSel}} != 3'b000));
  assign EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_valid = (EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_fire && EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD);
  assign EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_payload_robId = EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_fire = (EU0_ExecutionUnitBase_pipeline_execute_2_isFireing && ({EU0_CsrAccessPlugin_logic_wake_wakeRegFileSel,{EU0_DivPlugin_logic_wake_wakeRegFileSel,EU0_MulPlugin_logic_wake_wakeRegFileSel}} != 3'b000));
  assign EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_valid = (EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_fire && EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD);
  assign EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_payload_physical = EU0_ExecutionUnitBase_pipeline_execute_2_PHYS_RD;
  assign EU0_ExecutionUnitBase_pipeline_execute_2_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_execute_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_isRemoved = (EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed || EU0_ExecutionUnitBase_pipeline_execute_0_isThrown);
  assign EU0_ExecutionUnitBase_pipeline_execute_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_isThrown = 1'b0;
  assign EU0_ExecutionUnitBase_pipeline_fetch_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign EU0_ExecutionUnitBase_pipeline_fetch_0_ready = EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output;
  assign EU0_ExecutionUnitBase_pipeline_fetch_1_ready = EU0_ExecutionUnitBase_pipeline_fetch_1_ready_output;
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_1_valid = EU0_ExecutionUnitBase_pipeline_execute_0_valid;
    if(when_Pipeline_l278_2) begin
      _zz_EU0_ExecutionUnitBase_pipeline_execute_1_valid = 1'b0;
    end
  end

  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_0_ready = EU0_ExecutionUnitBase_pipeline_execute_0_ready_output;
    if(when_Pipeline_l278_2) begin
      EU0_ExecutionUnitBase_pipeline_execute_0_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_2 = (EU0_ExecutionUnitBase_pipeline_execute_0_haltRequest_DivPlugin_l83 != 1'b0);
  always @(*) begin
    _zz_EU0_ExecutionUnitBase_pipeline_execute_2_valid = EU0_ExecutionUnitBase_pipeline_execute_1_valid;
    if(when_Pipeline_l278_3) begin
      _zz_EU0_ExecutionUnitBase_pipeline_execute_2_valid = 1'b0;
    end
  end

  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_1_ready = EU0_ExecutionUnitBase_pipeline_execute_1_ready_output;
    if(when_Pipeline_l278_3) begin
      EU0_ExecutionUnitBase_pipeline_execute_1_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_3 = (EU0_ExecutionUnitBase_pipeline_execute_1_haltRequest_DivPlugin_l91 != 1'b0);
  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_2_ready = 1'b1;
    if(when_Pipeline_l278_4) begin
      EU0_ExecutionUnitBase_pipeline_execute_2_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_4 = ({EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_ExecutionUnitBase_l303,EU0_ExecutionUnitBase_pipeline_execute_2_haltRequest_CsrAccessPlugin_l373} != 2'b00);
  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output = EU0_ExecutionUnitBase_pipeline_fetch_1_ready;
    if(when_Connection_l74_1) begin
      EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_1 = (! EU0_ExecutionUnitBase_pipeline_fetch_1_valid);
  assign EU0_ExecutionUnitBase_pipeline_fetch_1_ready_output = EU0_ExecutionUnitBase_pipeline_execute_0_ready;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_valid = EU0_ExecutionUnitBase_pipeline_fetch_1_valid;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC2 = EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_REVERT = EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_ZERO = EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_SrcStageables_SRC1 = EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1 = EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS1;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS2 = EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS2;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS1_SIGNED = EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS1_SIGNED;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_RsUnsignedPlugin_RS2_SIGNED = EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS2_SIGNED;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM = EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_REM;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL = EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP = EU0_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SEL = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID = EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_ROB_MSB = EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_MSB;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_SC = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SC;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_AMO = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_AMO;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD = EU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD = EU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_LSU_ID = EU0_ExecutionUnitBase_pipeline_fetch_1_LSU_ID;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_PC = EU0_ExecutionUnitBase_pipeline_fetch_1_PC;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LR = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LR;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_AguPlugin_LOAD = EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LOAD;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_IMM = EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_IMM;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK = EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_MASK;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL = EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_CLEAR = EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_CLEAR;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_SEL = EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_SEL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_HIGH = EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_HIGH;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_EBREAK = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_EBREAK;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_ECALL = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_ECALL;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_XRET = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_XRET;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_I = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_I;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FLUSH_DATA = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FLUSH_DATA;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_VMA = EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_VMA;
  assign EU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E2 = EU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E2;
  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_0_ready_output = EU0_ExecutionUnitBase_pipeline_execute_1_ready;
    if(when_Connection_l74_2) begin
      EU0_ExecutionUnitBase_pipeline_execute_0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_2 = (! EU0_ExecutionUnitBase_pipeline_execute_1_valid);
  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_execute_1_ready_output = EU0_ExecutionUnitBase_pipeline_execute_2_ready;
    if(when_Connection_l74_3) begin
      EU0_ExecutionUnitBase_pipeline_execute_1_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_3 = (! EU0_ExecutionUnitBase_pipeline_execute_2_valid);
  assign BranchContextPlugin_free_dispatchMem_writes_0_port_valid = ((FrontendPlugin_dispatch_isFireing && FrontendPlugin_dispatch_BRANCH_SEL_0) && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0);
  assign BranchContextPlugin_free_dispatchMem_writes_0_port_payload_address = FrontendPlugin_dispatch_BRANCH_ID_0;
  assign BranchContextPlugin_free_dispatchMem_writes_0_port_payload_data = {FrontendPlugin_dispatch_Prediction_IS_BRANCH_0,{{FrontendPlugin_dispatch_GSHARE_COUNTER_0_1,FrontendPlugin_dispatch_GSHARE_COUNTER_0_0},FrontendPlugin_dispatch_BRANCH_HISTORY_0}};
  assign BranchContextPlugin_free_dispatchMem_writes_1_port_valid = ((FrontendPlugin_dispatch_isFireing && FrontendPlugin_dispatch_BRANCH_SEL_1) && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1);
  assign BranchContextPlugin_free_dispatchMem_writes_1_port_payload_address = FrontendPlugin_dispatch_BRANCH_ID_1;
  assign BranchContextPlugin_free_dispatchMem_writes_1_port_payload_data = {FrontendPlugin_dispatch_Prediction_IS_BRANCH_1,{{FrontendPlugin_dispatch_GSHARE_COUNTER_1_1,FrontendPlugin_dispatch_GSHARE_COUNTER_1_0},FrontendPlugin_dispatch_BRANCH_HISTORY_1}};
  assign BranchContextPlugin_free_learn_valid = (BranchContextPlugin_logic_ptr_free != BranchContextPlugin_logic_ptr_commited);
  assign BranchContextPlugin_free_learn_bid = BranchContextPlugin_logic_ptr_free[3:0];
  assign _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice = BranchContextPlugin_logic_mem_finalBranch_io_read_0_rsp;
  assign BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice = _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[31 : 0];
  assign BranchContextPlugin_learn_BRANCH_FINAL_pcTarget = _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[63 : 32];
  assign BranchContextPlugin_learn_BRANCH_FINAL_taken = _zz_BranchContextPlugin_learn_BRANCH_FINAL_pcOnLastSlice[64];
  assign BranchContextPlugin_free_learn_raw = BranchContextPlugin_free_dispatchMem_mem_io_read_0_rsp;
  assign BranchContextPlugin_free_learn_BRANCH_HISTORY = BranchContextPlugin_free_learn_raw[23 : 0];
  assign _zz_BranchContextPlugin_free_learn_GSHARE_COUNTER_0 = BranchContextPlugin_free_learn_raw[27 : 24];
  assign BranchContextPlugin_free_learn_GSHARE_COUNTER_0 = _zz_BranchContextPlugin_free_learn_GSHARE_COUNTER_0[1 : 0];
  assign BranchContextPlugin_free_learn_GSHARE_COUNTER_1 = _zz_BranchContextPlugin_free_learn_GSHARE_COUNTER_0[3 : 2];
  assign BranchContextPlugin_free_learn_Prediction_IS_BRANCH = BranchContextPlugin_free_learn_raw[28];
  assign BranchContextPlugin_setup_learnValid = BranchContextPlugin_free_learn_valid;
  assign DispatchPlugin_logic_queueStaticWakeTransposed_0 = {DispatchPlugin_logic_queue_io_contexts_31_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_30_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_29_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_28_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_27_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_26_staticWake[0],{DispatchPlugin_logic_queue_io_contexts_25_staticWake[0],{_zz_DispatchPlugin_logic_queueStaticWakeTransposed_0,{_zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_1,_zz_DispatchPlugin_logic_queueStaticWakeTransposed_0_2}}}}}}}}};
  assign DispatchPlugin_logic_queueStaticWakeTransposedHistory_0_0 = DispatchPlugin_logic_queueStaticWakeTransposed_0;
  assign toplevel_DispatchPlugin_logic_queue_io_push_fire = (FrontendPlugin_dispatch_isFireing && DispatchPlugin_logic_queue_io_push_ready);
  assign FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l187 = (! DispatchPlugin_logic_queue_io_push_ready);
  assign DispatchPlugin_logic_push_skip = (! ({FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1,FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0} != 2'b00));
  assign DispatchPlugin_logic_push_fenceOlder = (FrontendPlugin_dispatch_valid && ({(FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1 && FrontendPlugin_dispatch_DispatchPlugin_FENCE_OLDER_1),(FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 && FrontendPlugin_dispatch_DispatchPlugin_FENCE_OLDER_0)} != 2'b00));
  assign DispatchPlugin_logic_push_fenceYounger = (FrontendPlugin_dispatch_valid && ({(FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1 && FrontendPlugin_dispatch_DispatchPlugin_FENCE_YOUNGER_1),(FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 && FrontendPlugin_dispatch_DispatchPlugin_FENCE_YOUNGER_0)} != 2'b00));
  assign when_DispatchPlugin_l192 = (FrontendPlugin_dispatch_isFireing && (! DispatchPlugin_logic_push_skip));
  assign DispatchPlugin_logic_push_commitNotWaitingOnUs = (|_zz_DispatchPlugin_logic_push_commitNotWaitingOnUs);
  assign FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l195 = (DispatchPlugin_logic_push_fenceOlder && DispatchPlugin_logic_push_commitNotWaitingOnUs);
  assign FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l196 = ((DispatchPlugin_logic_push_fenceYoungerLast && DispatchPlugin_logic_push_commitNotWaitingOnUs) && (! DispatchPlugin_logic_push_skip));
  assign DispatchPlugin_logic_push_slots_0_self = ((FrontendPlugin_dispatch_WRITE_RD_0 && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) ? 32'h40000000 : 32'h00000000);
  assign DispatchPlugin_logic_push_slots_0_events_0 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_0 ? _zz_DispatchPlugin_logic_push_slots_0_events_0 : 32'h00000000);
  assign DispatchPlugin_logic_push_slots_0_events_1 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_0 ? _zz_DispatchPlugin_logic_push_slots_0_events_1 : 32'h00000000);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_0_event = ((DispatchPlugin_logic_push_slots_0_self | DispatchPlugin_logic_push_slots_0_events_0) | DispatchPlugin_logic_push_slots_0_events_1);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_0_sel = (FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 ? {FrontendPlugin_dispatch_EU0_SEL_0,FrontendPlugin_dispatch_ALU0_ALU1_SEL_0} : 2'b00);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_0_context_robId = (FrontendPlugin_dispatch_ROB_ID | 6'h00);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_0_context_staticWake[0] = (FrontendPlugin_dispatch_WRITE_RD_0 && FrontendPlugin_dispatch_LATENCY_0_0);
  assign DispatchPlugin_logic_push_slots_1_self = ((FrontendPlugin_dispatch_WRITE_RD_1 && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1) ? 32'h80000000 : 32'h00000000);
  assign DispatchPlugin_logic_push_slots_1_events_0 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_1 ? _zz_DispatchPlugin_logic_push_slots_1_events_0 : 32'h00000000);
  assign DispatchPlugin_logic_push_slots_1_events_1 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_1 ? _zz_DispatchPlugin_logic_push_slots_1_events_1 : 32'h00000000);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_1_event = ((DispatchPlugin_logic_push_slots_1_self | DispatchPlugin_logic_push_slots_1_events_0) | DispatchPlugin_logic_push_slots_1_events_1);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_1_sel = (FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1 ? {FrontendPlugin_dispatch_EU0_SEL_1,FrontendPlugin_dispatch_ALU0_ALU1_SEL_1} : 2'b00);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_1_context_robId = (FrontendPlugin_dispatch_ROB_ID | 6'h01);
  assign DispatchPlugin_logic_queue_io_push_payload_slots_1_context_staticWake[0] = (FrontendPlugin_dispatch_WRITE_RD_1 && FrontendPlugin_dispatch_LATENCY_0_1);
  assign DispatchPlugin_logic_pop_0_portEventFull = {1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[15],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[14],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[13],{1'b0,{DispatchPlugin_logic_queue_io_schedules_0_payload_event[12],{_zz_DispatchPlugin_logic_pop_0_portEventFull,{_zz_DispatchPlugin_logic_pop_0_portEventFull_1,_zz_DispatchPlugin_logic_pop_0_portEventFull_2}}}}}}}}}};
  assign DispatchPlugin_logic_pop_0_stagesList_0_valid = DispatchPlugin_logic_queue_io_schedules_0_valid;
  assign DispatchPlugin_logic_pop_0_stagesList_0_OH = DispatchPlugin_logic_pop_0_portEventFull;
  assign DispatchPlugin_logic_pop_0_stagesList_0_OFFSET = DispatchPlugin_logic_ptr_current;
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT = DispatchPlugin_logic_pop_0_stagesList_0_OH[3];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_1 = DispatchPlugin_logic_pop_0_stagesList_0_OH[5];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_2 = DispatchPlugin_logic_pop_0_stagesList_0_OH[6];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3 = DispatchPlugin_logic_pop_0_stagesList_0_OH[7];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_4 = DispatchPlugin_logic_pop_0_stagesList_0_OH[9];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_5 = DispatchPlugin_logic_pop_0_stagesList_0_OH[10];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_6 = DispatchPlugin_logic_pop_0_stagesList_0_OH[11];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_7 = DispatchPlugin_logic_pop_0_stagesList_0_OH[12];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_8 = DispatchPlugin_logic_pop_0_stagesList_0_OH[13];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_9 = DispatchPlugin_logic_pop_0_stagesList_0_OH[14];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_10 = DispatchPlugin_logic_pop_0_stagesList_0_OH[15];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_11 = DispatchPlugin_logic_pop_0_stagesList_0_OH[17];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_12 = DispatchPlugin_logic_pop_0_stagesList_0_OH[18];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_13 = DispatchPlugin_logic_pop_0_stagesList_0_OH[19];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_14 = DispatchPlugin_logic_pop_0_stagesList_0_OH[20];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_15 = DispatchPlugin_logic_pop_0_stagesList_0_OH[21];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_16 = DispatchPlugin_logic_pop_0_stagesList_0_OH[22];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_17 = DispatchPlugin_logic_pop_0_stagesList_0_OH[23];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_18 = DispatchPlugin_logic_pop_0_stagesList_0_OH[24];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_19 = DispatchPlugin_logic_pop_0_stagesList_0_OH[25];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_20 = DispatchPlugin_logic_pop_0_stagesList_0_OH[26];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_21 = DispatchPlugin_logic_pop_0_stagesList_0_OH[27];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_22 = DispatchPlugin_logic_pop_0_stagesList_0_OH[28];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_23 = DispatchPlugin_logic_pop_0_stagesList_0_OH[29];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_24 = DispatchPlugin_logic_pop_0_stagesList_0_OH[30];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_25 = DispatchPlugin_logic_pop_0_stagesList_0_OH[31];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_26 = (((((((((((((((DispatchPlugin_logic_pop_0_stagesList_0_OH[1] || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_4) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_6) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_8) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_11) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_13) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_15) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_19) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_27 = (((((((((((((((DispatchPlugin_logic_pop_0_stagesList_0_OH[2] || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_5) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_6) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_9) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_12) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_13) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_16) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_20) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_28 = (((((((((((((((DispatchPlugin_logic_pop_0_stagesList_0_OH[4] || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_3) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_7) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_8) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_9) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_14) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_15) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_16) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_22) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_29 = (((((((((((((((DispatchPlugin_logic_pop_0_stagesList_0_OH[8] || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_4) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_5) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_6) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_7) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_8) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_9) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_18) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_19) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_20) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_22) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_30 = (((((((((((((((DispatchPlugin_logic_pop_0_stagesList_0_OH[16] || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_11) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_12) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_13) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_14) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_15) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_16) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_18) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_19) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_20) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_22) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_25);
  assign DispatchPlugin_logic_pop_0_stagesList_0_UINT = {_zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_30,{_zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_29,{_zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_28,{_zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_27,_zz_DispatchPlugin_logic_pop_0_stagesList_0_UINT_26}}}};
  assign DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID = (_zz_DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID + DispatchPlugin_logic_pop_0_stagesList_1_OFFSET);
  assign DispatchPlugin_logic_pop_0_stagesList_0_LATENCY_0 = (|(DispatchPlugin_logic_pop_0_stagesList_0_OH & DispatchPlugin_logic_queueStaticWakeTransposedHistory_0_0));
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[2 : 0];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[5 : 3];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[8 : 6];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[11 : 9];
  assign _zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_4 = DispatchPlugin_logic_queue_io_schedules_0_payload_event[14 : 12];
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0 = (((_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0[0] ? DispatchPlugin_logic_queue_io_contexts_0_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0[1] ? DispatchPlugin_logic_queue_io_contexts_2_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0[2] ? DispatchPlugin_logic_queue_io_contexts_4_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1 = (((_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1[0] ? DispatchPlugin_logic_queue_io_contexts_6_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1[1] ? DispatchPlugin_logic_queue_io_contexts_8_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1[2] ? DispatchPlugin_logic_queue_io_contexts_10_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2 = (((_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2[0] ? DispatchPlugin_logic_queue_io_contexts_12_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2[1] ? DispatchPlugin_logic_queue_io_contexts_14_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2[2] ? DispatchPlugin_logic_queue_io_contexts_16_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3 = (((_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3[0] ? DispatchPlugin_logic_queue_io_contexts_18_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3[1] ? DispatchPlugin_logic_queue_io_contexts_20_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3[2] ? DispatchPlugin_logic_queue_io_contexts_22_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_4 = (((_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_4[0] ? DispatchPlugin_logic_queue_io_contexts_24_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_4[1] ? DispatchPlugin_logic_queue_io_contexts_26_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_4[2] ? DispatchPlugin_logic_queue_io_contexts_28_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_5 = (DispatchPlugin_logic_queue_io_schedules_0_payload_event[15] ? DispatchPlugin_logic_queue_io_contexts_30_physRd : 6'h00);
  assign DispatchPlugin_logic_pop_0_stagesList_1_PHYS_RD = (((DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_0 | DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_1) | (DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_2 | DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_3)) | (DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_4 | DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_5));
  assign ALU0_ExecutionUnitBase_pipeline_push_port_valid = DispatchPlugin_logic_pop_0_stagesList_1_valid;
  assign ALU0_ExecutionUnitBase_pipeline_push_port_robId = DispatchPlugin_logic_pop_0_stagesList_1_ROB_ID;
  assign ALU0_ExecutionUnitBase_pipeline_push_port_physRd = DispatchPlugin_logic_pop_0_stagesList_1_PHYS_RD;
  assign toplevel_DispatchPlugin_logic_queue_io_schedules_0_fire = (DispatchPlugin_logic_queue_io_schedules_0_valid && DispatchPlugin_logic_pop_0_stagesList_0_ready);
  assign DispatchPlugin_logic_pop_0_wake_L0_mask = (toplevel_DispatchPlugin_logic_queue_io_schedules_0_fire ? DispatchPlugin_logic_pop_0_portEventFull : 32'h00000000);
  assign DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid = (DispatchPlugin_logic_pop_0_stagesList_1_valid && DispatchPlugin_logic_pop_0_stagesList_1_LATENCY_0);
  assign DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical = DispatchPlugin_logic_pop_0_stagesList_1_PHYS_RD;
  assign DispatchPlugin_logic_pop_0_stagesList_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_0_stagesList_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_0_stagesList_0_ready = 1'b1;
  assign DispatchPlugin_logic_pop_1_portEventFull = {DispatchPlugin_logic_queue_io_schedules_1_payload_event[15],{1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[14],{1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[13],{1'b0,{DispatchPlugin_logic_queue_io_schedules_1_payload_event[12],{1'b0,{_zz_DispatchPlugin_logic_pop_1_portEventFull,{_zz_DispatchPlugin_logic_pop_1_portEventFull_1,_zz_DispatchPlugin_logic_pop_1_portEventFull_2}}}}}}}}}};
  assign DispatchPlugin_logic_pop_1_stagesList_0_valid = DispatchPlugin_logic_queue_io_schedules_1_valid;
  assign DispatchPlugin_logic_pop_1_stagesList_0_OH = DispatchPlugin_logic_pop_1_portEventFull;
  assign DispatchPlugin_logic_pop_1_stagesList_0_OFFSET = DispatchPlugin_logic_ptr_current;
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT = DispatchPlugin_logic_pop_1_stagesList_0_OH[3];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_1 = DispatchPlugin_logic_pop_1_stagesList_0_OH[5];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_2 = DispatchPlugin_logic_pop_1_stagesList_0_OH[6];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3 = DispatchPlugin_logic_pop_1_stagesList_0_OH[7];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_4 = DispatchPlugin_logic_pop_1_stagesList_0_OH[9];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_5 = DispatchPlugin_logic_pop_1_stagesList_0_OH[10];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_6 = DispatchPlugin_logic_pop_1_stagesList_0_OH[11];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_7 = DispatchPlugin_logic_pop_1_stagesList_0_OH[12];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_8 = DispatchPlugin_logic_pop_1_stagesList_0_OH[13];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_9 = DispatchPlugin_logic_pop_1_stagesList_0_OH[14];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_10 = DispatchPlugin_logic_pop_1_stagesList_0_OH[15];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_11 = DispatchPlugin_logic_pop_1_stagesList_0_OH[17];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_12 = DispatchPlugin_logic_pop_1_stagesList_0_OH[18];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_13 = DispatchPlugin_logic_pop_1_stagesList_0_OH[19];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_14 = DispatchPlugin_logic_pop_1_stagesList_0_OH[20];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_15 = DispatchPlugin_logic_pop_1_stagesList_0_OH[21];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_16 = DispatchPlugin_logic_pop_1_stagesList_0_OH[22];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_17 = DispatchPlugin_logic_pop_1_stagesList_0_OH[23];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_18 = DispatchPlugin_logic_pop_1_stagesList_0_OH[24];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_19 = DispatchPlugin_logic_pop_1_stagesList_0_OH[25];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_20 = DispatchPlugin_logic_pop_1_stagesList_0_OH[26];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_21 = DispatchPlugin_logic_pop_1_stagesList_0_OH[27];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_22 = DispatchPlugin_logic_pop_1_stagesList_0_OH[28];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_23 = DispatchPlugin_logic_pop_1_stagesList_0_OH[29];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_24 = DispatchPlugin_logic_pop_1_stagesList_0_OH[30];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_25 = DispatchPlugin_logic_pop_1_stagesList_0_OH[31];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_26 = (((((((((((((((DispatchPlugin_logic_pop_1_stagesList_0_OH[1] || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_4) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_6) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_8) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_11) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_13) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_15) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_19) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_27 = (((((((((((((((DispatchPlugin_logic_pop_1_stagesList_0_OH[2] || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_5) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_6) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_9) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_12) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_13) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_16) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_20) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_28 = (((((((((((((((DispatchPlugin_logic_pop_1_stagesList_0_OH[4] || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_3) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_7) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_8) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_9) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_14) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_15) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_16) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_22) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_29 = (((((((((((((((DispatchPlugin_logic_pop_1_stagesList_0_OH[8] || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_4) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_5) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_6) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_7) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_8) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_9) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_18) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_19) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_20) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_22) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_30 = (((((((((((((((DispatchPlugin_logic_pop_1_stagesList_0_OH[16] || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_11) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_12) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_13) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_14) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_15) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_16) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_18) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_19) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_20) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_22) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_25);
  assign DispatchPlugin_logic_pop_1_stagesList_0_UINT = {_zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_30,{_zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_29,{_zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_28,{_zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_27,_zz_DispatchPlugin_logic_pop_1_stagesList_0_UINT_26}}}};
  assign DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID = (_zz_DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID + DispatchPlugin_logic_pop_1_stagesList_1_OFFSET);
  assign DispatchPlugin_logic_pop_1_stagesList_0_LATENCY_0 = (|(DispatchPlugin_logic_pop_1_stagesList_0_OH & DispatchPlugin_logic_queueStaticWakeTransposedHistory_0_0));
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_0 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[2 : 0];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_1 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[5 : 3];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_2 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[8 : 6];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_3 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[11 : 9];
  assign _zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_4 = DispatchPlugin_logic_queue_io_schedules_1_payload_event[14 : 12];
  assign DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_0 = (((_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_0[0] ? DispatchPlugin_logic_queue_io_contexts_1_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_0[1] ? DispatchPlugin_logic_queue_io_contexts_3_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_0[2] ? DispatchPlugin_logic_queue_io_contexts_5_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_1 = (((_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_1[0] ? DispatchPlugin_logic_queue_io_contexts_7_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_1[1] ? DispatchPlugin_logic_queue_io_contexts_9_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_1[2] ? DispatchPlugin_logic_queue_io_contexts_11_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_2 = (((_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_2[0] ? DispatchPlugin_logic_queue_io_contexts_13_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_2[1] ? DispatchPlugin_logic_queue_io_contexts_15_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_2[2] ? DispatchPlugin_logic_queue_io_contexts_17_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_3 = (((_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_3[0] ? DispatchPlugin_logic_queue_io_contexts_19_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_3[1] ? DispatchPlugin_logic_queue_io_contexts_21_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_3[2] ? DispatchPlugin_logic_queue_io_contexts_23_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_4 = (((_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_4[0] ? DispatchPlugin_logic_queue_io_contexts_25_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_4[1] ? DispatchPlugin_logic_queue_io_contexts_27_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_4[2] ? DispatchPlugin_logic_queue_io_contexts_29_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_5 = (DispatchPlugin_logic_queue_io_schedules_1_payload_event[15] ? DispatchPlugin_logic_queue_io_contexts_31_physRd : 6'h00);
  assign DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RD = (((DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_0 | DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_1) | (DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_2 | DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_3)) | (DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_4 | DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_5));
  assign ALU1_ExecutionUnitBase_pipeline_push_port_valid = DispatchPlugin_logic_pop_1_stagesList_1_valid;
  assign ALU1_ExecutionUnitBase_pipeline_push_port_robId = DispatchPlugin_logic_pop_1_stagesList_1_ROB_ID;
  assign ALU1_ExecutionUnitBase_pipeline_push_port_physRd = DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RD;
  assign toplevel_DispatchPlugin_logic_queue_io_schedules_1_fire = (DispatchPlugin_logic_queue_io_schedules_1_valid && DispatchPlugin_logic_pop_1_stagesList_0_ready);
  assign DispatchPlugin_logic_pop_1_wake_L0_mask = (toplevel_DispatchPlugin_logic_queue_io_schedules_1_fire ? DispatchPlugin_logic_pop_1_portEventFull : 32'h00000000);
  assign DispatchPlugin_logic_pop_1_wake_L0_bypassed_valid = (DispatchPlugin_logic_pop_1_stagesList_1_valid && DispatchPlugin_logic_pop_1_stagesList_1_LATENCY_0);
  assign DispatchPlugin_logic_pop_1_wake_L0_bypassed_payload_physical = DispatchPlugin_logic_pop_1_stagesList_1_PHYS_RD;
  assign DispatchPlugin_logic_pop_1_stagesList_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_1_stagesList_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_1_stagesList_0_ready = 1'b1;
  assign DispatchPlugin_logic_pop_2_portEventFull = {DispatchPlugin_logic_queue_io_schedules_2_payload_event[31],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[30],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[29],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[28],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[27],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[26],{DispatchPlugin_logic_queue_io_schedules_2_payload_event[25],{_zz_DispatchPlugin_logic_pop_2_portEventFull,{_zz_DispatchPlugin_logic_pop_2_portEventFull_1,_zz_DispatchPlugin_logic_pop_2_portEventFull_2}}}}}}}}};
  assign DispatchPlugin_logic_pop_2_stagesList_0_valid = DispatchPlugin_logic_queue_io_schedules_2_valid;
  assign DispatchPlugin_logic_pop_2_stagesList_0_OH = DispatchPlugin_logic_pop_2_portEventFull;
  assign DispatchPlugin_logic_pop_2_stagesList_0_OFFSET = DispatchPlugin_logic_ptr_current;
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT = DispatchPlugin_logic_pop_2_stagesList_0_OH[3];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_1 = DispatchPlugin_logic_pop_2_stagesList_0_OH[5];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_2 = DispatchPlugin_logic_pop_2_stagesList_0_OH[6];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_3 = DispatchPlugin_logic_pop_2_stagesList_0_OH[7];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_4 = DispatchPlugin_logic_pop_2_stagesList_0_OH[9];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_5 = DispatchPlugin_logic_pop_2_stagesList_0_OH[10];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_6 = DispatchPlugin_logic_pop_2_stagesList_0_OH[11];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_7 = DispatchPlugin_logic_pop_2_stagesList_0_OH[12];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_8 = DispatchPlugin_logic_pop_2_stagesList_0_OH[13];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_9 = DispatchPlugin_logic_pop_2_stagesList_0_OH[14];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_10 = DispatchPlugin_logic_pop_2_stagesList_0_OH[15];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_11 = DispatchPlugin_logic_pop_2_stagesList_0_OH[17];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_12 = DispatchPlugin_logic_pop_2_stagesList_0_OH[18];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_13 = DispatchPlugin_logic_pop_2_stagesList_0_OH[19];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_14 = DispatchPlugin_logic_pop_2_stagesList_0_OH[20];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_15 = DispatchPlugin_logic_pop_2_stagesList_0_OH[21];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_16 = DispatchPlugin_logic_pop_2_stagesList_0_OH[22];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_17 = DispatchPlugin_logic_pop_2_stagesList_0_OH[23];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_18 = DispatchPlugin_logic_pop_2_stagesList_0_OH[24];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_19 = DispatchPlugin_logic_pop_2_stagesList_0_OH[25];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_20 = DispatchPlugin_logic_pop_2_stagesList_0_OH[26];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_21 = DispatchPlugin_logic_pop_2_stagesList_0_OH[27];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_22 = DispatchPlugin_logic_pop_2_stagesList_0_OH[28];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_23 = DispatchPlugin_logic_pop_2_stagesList_0_OH[29];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_24 = DispatchPlugin_logic_pop_2_stagesList_0_OH[30];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_25 = DispatchPlugin_logic_pop_2_stagesList_0_OH[31];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_26 = (((((((((((((((DispatchPlugin_logic_pop_2_stagesList_0_OH[1] || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_3) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_4) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_6) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_8) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_11) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_13) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_15) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_19) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_27 = (((((((((((((((DispatchPlugin_logic_pop_2_stagesList_0_OH[2] || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_3) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_5) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_6) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_9) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_12) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_13) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_16) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_20) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_28 = (((((((((((((((DispatchPlugin_logic_pop_2_stagesList_0_OH[4] || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_1) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_2) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_3) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_7) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_8) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_9) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_14) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_15) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_16) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_22) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_29 = (((((((((((((((DispatchPlugin_logic_pop_2_stagesList_0_OH[8] || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_4) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_5) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_6) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_7) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_8) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_9) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_10) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_18) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_19) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_20) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_22) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_25);
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_30 = (((((((((((((((DispatchPlugin_logic_pop_2_stagesList_0_OH[16] || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_11) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_12) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_13) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_14) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_15) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_16) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_17) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_18) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_19) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_20) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_21) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_22) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_23) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_24) || _zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_25);
  assign DispatchPlugin_logic_pop_2_stagesList_0_UINT = {_zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_30,{_zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_29,{_zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_28,{_zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_27,_zz_DispatchPlugin_logic_pop_2_stagesList_0_UINT_26}}}};
  assign DispatchPlugin_logic_pop_2_stagesList_1_ROB_ID = (_zz_DispatchPlugin_logic_pop_2_stagesList_1_ROB_ID + DispatchPlugin_logic_pop_2_stagesList_1_OFFSET);
  assign DispatchPlugin_logic_pop_2_stagesList_0_LATENCY_0 = (|(DispatchPlugin_logic_pop_2_stagesList_0_OH & DispatchPlugin_logic_queueStaticWakeTransposedHistory_0_0));
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_0 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[2 : 0];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_1 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[5 : 3];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_2 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[8 : 6];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_3 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[11 : 9];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_4 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[14 : 12];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_5 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[17 : 15];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_6 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[20 : 18];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_7 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[23 : 21];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_8 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[26 : 24];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_9 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[29 : 27];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_10 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[31 : 30];
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_0 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_0[0] ? DispatchPlugin_logic_queue_io_contexts_0_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_0[1] ? DispatchPlugin_logic_queue_io_contexts_1_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_0[2] ? DispatchPlugin_logic_queue_io_contexts_2_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_1 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_1[0] ? DispatchPlugin_logic_queue_io_contexts_3_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_1[1] ? DispatchPlugin_logic_queue_io_contexts_4_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_1[2] ? DispatchPlugin_logic_queue_io_contexts_5_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_2 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_2[0] ? DispatchPlugin_logic_queue_io_contexts_6_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_2[1] ? DispatchPlugin_logic_queue_io_contexts_7_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_2[2] ? DispatchPlugin_logic_queue_io_contexts_8_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_3 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_3[0] ? DispatchPlugin_logic_queue_io_contexts_9_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_3[1] ? DispatchPlugin_logic_queue_io_contexts_10_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_3[2] ? DispatchPlugin_logic_queue_io_contexts_11_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_4 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_4[0] ? DispatchPlugin_logic_queue_io_contexts_12_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_4[1] ? DispatchPlugin_logic_queue_io_contexts_13_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_4[2] ? DispatchPlugin_logic_queue_io_contexts_14_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_5 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_5[0] ? DispatchPlugin_logic_queue_io_contexts_15_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_5[1] ? DispatchPlugin_logic_queue_io_contexts_16_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_5[2] ? DispatchPlugin_logic_queue_io_contexts_17_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_6 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_6[0] ? DispatchPlugin_logic_queue_io_contexts_18_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_6[1] ? DispatchPlugin_logic_queue_io_contexts_19_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_6[2] ? DispatchPlugin_logic_queue_io_contexts_20_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_7 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_7[0] ? DispatchPlugin_logic_queue_io_contexts_21_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_7[1] ? DispatchPlugin_logic_queue_io_contexts_22_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_7[2] ? DispatchPlugin_logic_queue_io_contexts_23_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_8 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_8[0] ? DispatchPlugin_logic_queue_io_contexts_24_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_8[1] ? DispatchPlugin_logic_queue_io_contexts_25_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_8[2] ? DispatchPlugin_logic_queue_io_contexts_26_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_9 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_9[0] ? DispatchPlugin_logic_queue_io_contexts_27_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_9[1] ? DispatchPlugin_logic_queue_io_contexts_28_physRd : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_9[2] ? DispatchPlugin_logic_queue_io_contexts_29_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_10 = ((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_10[0] ? DispatchPlugin_logic_queue_io_contexts_30_physRd : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_10[1] ? DispatchPlugin_logic_queue_io_contexts_31_physRd : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_1_PHYS_RD = ((((DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_0 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_1) | (DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_2 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_3)) | ((DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_4 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_5) | (DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_6 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_7))) | ((DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_8 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_9) | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_10));
  assign EU0_ExecutionUnitBase_pipeline_push_port_valid = DispatchPlugin_logic_pop_2_stagesList_1_valid;
  assign EU0_ExecutionUnitBase_pipeline_push_port_robId = DispatchPlugin_logic_pop_2_stagesList_1_ROB_ID;
  assign EU0_ExecutionUnitBase_pipeline_push_port_physRd = DispatchPlugin_logic_pop_2_stagesList_1_PHYS_RD;
  assign DispatchPlugin_logic_pop_2_stagesList_1_haltRequest_DispatchPlugin_l292 = (! EU0_ExecutionUnitBase_pipeline_push_port_ready);
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_0 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[2 : 0];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_1 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[5 : 3];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_2 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[8 : 6];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_3 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[11 : 9];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_4 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[14 : 12];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_5 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[17 : 15];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_6 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[20 : 18];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_7 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[23 : 21];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_8 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[26 : 24];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_9 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[29 : 27];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_10 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[31 : 30];
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_0 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_0[0] ? DispatchPlugin_logic_queue_io_contexts_0_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_0[1] ? DispatchPlugin_logic_queue_io_contexts_1_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_0[2] ? DispatchPlugin_logic_queue_io_contexts_2_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_1 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_1[0] ? DispatchPlugin_logic_queue_io_contexts_3_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_1[1] ? DispatchPlugin_logic_queue_io_contexts_4_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_1[2] ? DispatchPlugin_logic_queue_io_contexts_5_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_2 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_2[0] ? DispatchPlugin_logic_queue_io_contexts_6_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_2[1] ? DispatchPlugin_logic_queue_io_contexts_7_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_2[2] ? DispatchPlugin_logic_queue_io_contexts_8_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_3 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_3[0] ? DispatchPlugin_logic_queue_io_contexts_9_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_3[1] ? DispatchPlugin_logic_queue_io_contexts_10_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_3[2] ? DispatchPlugin_logic_queue_io_contexts_11_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_4 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_4[0] ? DispatchPlugin_logic_queue_io_contexts_12_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_4[1] ? DispatchPlugin_logic_queue_io_contexts_13_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_4[2] ? DispatchPlugin_logic_queue_io_contexts_14_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_5 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_5[0] ? DispatchPlugin_logic_queue_io_contexts_15_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_5[1] ? DispatchPlugin_logic_queue_io_contexts_16_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_5[2] ? DispatchPlugin_logic_queue_io_contexts_17_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_6 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_6[0] ? DispatchPlugin_logic_queue_io_contexts_18_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_6[1] ? DispatchPlugin_logic_queue_io_contexts_19_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_6[2] ? DispatchPlugin_logic_queue_io_contexts_20_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_7 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_7[0] ? DispatchPlugin_logic_queue_io_contexts_21_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_7[1] ? DispatchPlugin_logic_queue_io_contexts_22_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_7[2] ? DispatchPlugin_logic_queue_io_contexts_23_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_8 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_8[0] ? DispatchPlugin_logic_queue_io_contexts_24_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_8[1] ? DispatchPlugin_logic_queue_io_contexts_25_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_8[2] ? DispatchPlugin_logic_queue_io_contexts_26_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_9 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_9[0] ? DispatchPlugin_logic_queue_io_contexts_27_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_9[1] ? DispatchPlugin_logic_queue_io_contexts_28_euCtx_0 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_9[2] ? DispatchPlugin_logic_queue_io_contexts_29_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_10 = ((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_10[0] ? DispatchPlugin_logic_queue_io_contexts_30_euCtx_0 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_10[1] ? DispatchPlugin_logic_queue_io_contexts_31_euCtx_0 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_1_PHYS_RS_0 = ((((DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_0 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_1) | (DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_2 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_3)) | ((DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_4 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_5) | (DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_6 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_7))) | ((DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_8 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_9) | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_10));
  assign EU0_ExecutionUnitBase_pipeline_push_port_context_0 = DispatchPlugin_logic_pop_2_stagesList_1_PHYS_RS_0;
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_0 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[2 : 0];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_1 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[5 : 3];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_2 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[8 : 6];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_3 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[11 : 9];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_4 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[14 : 12];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_5 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[17 : 15];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_6 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[20 : 18];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_7 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[23 : 21];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_8 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[26 : 24];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_9 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[29 : 27];
  assign _zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_10 = DispatchPlugin_logic_queue_io_schedules_2_payload_event[31 : 30];
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_0 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_0[0] ? DispatchPlugin_logic_queue_io_contexts_0_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_0[1] ? DispatchPlugin_logic_queue_io_contexts_1_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_0[2] ? DispatchPlugin_logic_queue_io_contexts_2_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_1 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_1[0] ? DispatchPlugin_logic_queue_io_contexts_3_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_1[1] ? DispatchPlugin_logic_queue_io_contexts_4_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_1[2] ? DispatchPlugin_logic_queue_io_contexts_5_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_2 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_2[0] ? DispatchPlugin_logic_queue_io_contexts_6_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_2[1] ? DispatchPlugin_logic_queue_io_contexts_7_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_2[2] ? DispatchPlugin_logic_queue_io_contexts_8_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_3 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_3[0] ? DispatchPlugin_logic_queue_io_contexts_9_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_3[1] ? DispatchPlugin_logic_queue_io_contexts_10_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_3[2] ? DispatchPlugin_logic_queue_io_contexts_11_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_4 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_4[0] ? DispatchPlugin_logic_queue_io_contexts_12_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_4[1] ? DispatchPlugin_logic_queue_io_contexts_13_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_4[2] ? DispatchPlugin_logic_queue_io_contexts_14_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_5 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_5[0] ? DispatchPlugin_logic_queue_io_contexts_15_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_5[1] ? DispatchPlugin_logic_queue_io_contexts_16_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_5[2] ? DispatchPlugin_logic_queue_io_contexts_17_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_6 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_6[0] ? DispatchPlugin_logic_queue_io_contexts_18_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_6[1] ? DispatchPlugin_logic_queue_io_contexts_19_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_6[2] ? DispatchPlugin_logic_queue_io_contexts_20_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_7 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_7[0] ? DispatchPlugin_logic_queue_io_contexts_21_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_7[1] ? DispatchPlugin_logic_queue_io_contexts_22_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_7[2] ? DispatchPlugin_logic_queue_io_contexts_23_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_8 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_8[0] ? DispatchPlugin_logic_queue_io_contexts_24_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_8[1] ? DispatchPlugin_logic_queue_io_contexts_25_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_8[2] ? DispatchPlugin_logic_queue_io_contexts_26_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_9 = (((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_9[0] ? DispatchPlugin_logic_queue_io_contexts_27_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_9[1] ? DispatchPlugin_logic_queue_io_contexts_28_euCtx_1 : 6'h00)) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_9[2] ? DispatchPlugin_logic_queue_io_contexts_29_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_10 = ((_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_10[0] ? DispatchPlugin_logic_queue_io_contexts_30_euCtx_1 : 6'h00) | (_zz_DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_10[1] ? DispatchPlugin_logic_queue_io_contexts_31_euCtx_1 : 6'h00));
  assign DispatchPlugin_logic_pop_2_stagesList_1_PHYS_RS_1 = ((((DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_0 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_1) | (DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_2 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_3)) | ((DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_4 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_5) | (DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_6 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_7))) | ((DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_8 | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_9) | DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_10));
  assign EU0_ExecutionUnitBase_pipeline_push_port_context_1 = DispatchPlugin_logic_pop_2_stagesList_1_PHYS_RS_1;
  assign DispatchPlugin_logic_pop_2_stagesList_1_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_2_stagesList_0_isFlushed = CommitPlugin_logic_commit_reschedulePort_valid;
  assign DispatchPlugin_logic_pop_2_stagesList_0_ready = DispatchPlugin_logic_pop_2_stagesList_0_ready_output;
  always @(*) begin
    DispatchPlugin_logic_pop_2_stagesList_1_ready = 1'b1;
    if(when_Pipeline_l278_5) begin
      DispatchPlugin_logic_pop_2_stagesList_1_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_5 = (DispatchPlugin_logic_pop_2_stagesList_1_haltRequest_DispatchPlugin_l292 != 1'b0);
  always @(*) begin
    DispatchPlugin_logic_pop_2_stagesList_0_ready_output = DispatchPlugin_logic_pop_2_stagesList_1_ready;
    if(when_Connection_l74_4) begin
      DispatchPlugin_logic_pop_2_stagesList_0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_4 = (! DispatchPlugin_logic_pop_2_stagesList_1_valid);
  assign DispatchPlugin_logic_wake_dynamic_offseted_0_valid = Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRob_valid;
  assign DispatchPlugin_logic_wake_dynamic_offseted_0_payload = _zz_DispatchPlugin_logic_wake_dynamic_offseted_0_payload[4:0];
  assign DispatchPlugin_logic_wake_dynamic_offseted_1_valid = Lsu2Plugin_logic_sharedPip_ctrl_wakeRob_valid;
  assign DispatchPlugin_logic_wake_dynamic_offseted_1_payload = _zz_DispatchPlugin_logic_wake_dynamic_offseted_1_payload[4:0];
  assign DispatchPlugin_logic_wake_dynamic_offseted_2_valid = Lsu2Plugin_logic_special_wakeRob_valid;
  assign DispatchPlugin_logic_wake_dynamic_offseted_2_payload = _zz_DispatchPlugin_logic_wake_dynamic_offseted_2_payload[4:0];
  assign DispatchPlugin_logic_wake_dynamic_offseted_3_valid = EU0_ExecutionUnitBase_pipeline_wakeRobs_logic_0_rob_valid;
  assign DispatchPlugin_logic_wake_dynamic_offseted_3_payload = _zz_DispatchPlugin_logic_wake_dynamic_offseted_3_payload[4:0];
  assign DispatchPlugin_logic_wake_dynamic_masks_0 = ((DispatchPlugin_logic_wake_dynamic_offseted_0_valid ? 32'hffffffff : 32'h00000000) & _zz_DispatchPlugin_logic_wake_dynamic_masks_0);
  assign DispatchPlugin_logic_wake_dynamic_masks_1 = ((DispatchPlugin_logic_wake_dynamic_offseted_1_valid ? 32'hffffffff : 32'h00000000) & _zz_DispatchPlugin_logic_wake_dynamic_masks_1);
  assign DispatchPlugin_logic_wake_dynamic_masks_2 = ((DispatchPlugin_logic_wake_dynamic_offseted_2_valid ? 32'hffffffff : 32'h00000000) & _zz_DispatchPlugin_logic_wake_dynamic_masks_2);
  assign DispatchPlugin_logic_wake_dynamic_masks_3 = ((DispatchPlugin_logic_wake_dynamic_offseted_3_valid ? 32'hffffffff : 32'h00000000) & _zz_DispatchPlugin_logic_wake_dynamic_masks_3);
  assign DispatchPlugin_logic_wake_statics_0_popMask = ((DispatchPlugin_logic_pop_0_wake_L0_mask | DispatchPlugin_logic_pop_1_wake_L0_mask) & DispatchPlugin_logic_queueStaticWakeTransposed_0);
  assign DispatchPlugin_logic_wake_statics_0_history_0 = DispatchPlugin_logic_wake_statics_0_popMask;
  assign DispatchPlugin_logic_wake_optReduce_relaxed = ((DispatchPlugin_logic_wake_dynamic_masks_0 | DispatchPlugin_logic_wake_dynamic_masks_1) | (DispatchPlugin_logic_wake_dynamic_masks_2 | DispatchPlugin_logic_wake_dynamic_masks_3));
  assign DispatchPlugin_logic_wake_optReduce_reduced = (DispatchPlugin_logic_wake_optReduce_relaxed | DispatchPlugin_logic_wake_statics_0_history_0);
  assign DispatchPlugin_logic_whitebox_issuePorts_0_valid = (ALU0_ExecutionUnitBase_pipeline_push_port_valid && 1'b1);
  assign DispatchPlugin_logic_whitebox_issuePorts_0_payload_robId = ALU0_ExecutionUnitBase_pipeline_push_port_robId;
  assign DispatchPlugin_logic_whitebox_issuePorts_0_payload_physRd = ALU0_ExecutionUnitBase_pipeline_push_port_physRd;
  assign DispatchPlugin_logic_whitebox_issuePorts_1_valid = (ALU1_ExecutionUnitBase_pipeline_push_port_valid && 1'b1);
  assign DispatchPlugin_logic_whitebox_issuePorts_1_payload_robId = ALU1_ExecutionUnitBase_pipeline_push_port_robId;
  assign DispatchPlugin_logic_whitebox_issuePorts_1_payload_physRd = ALU1_ExecutionUnitBase_pipeline_push_port_physRd;
  assign DispatchPlugin_logic_whitebox_issuePorts_2_valid = (EU0_ExecutionUnitBase_pipeline_push_port_valid && EU0_ExecutionUnitBase_pipeline_push_port_ready);
  assign DispatchPlugin_logic_whitebox_issuePorts_2_payload_robId = EU0_ExecutionUnitBase_pipeline_push_port_robId;
  assign DispatchPlugin_logic_whitebox_issuePorts_2_payload_physRd = EU0_ExecutionUnitBase_pipeline_push_port_physRd;
  assign DispatchPlugin_logic_whitebox_issuePorts_2_payload_context_0 = EU0_ExecutionUnitBase_pipeline_push_port_context_0;
  assign DispatchPlugin_logic_whitebox_issuePorts_2_payload_context_1 = EU0_ExecutionUnitBase_pipeline_push_port_context_1;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_valid = (Lsu2Plugin_setup_regfilePorts_0_write_valid != 1'b0);
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_address = Lsu2Plugin_setup_regfilePorts_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_data = Lsu2Plugin_setup_regfilePorts_0_write_data;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_robId = Lsu2Plugin_setup_regfilePorts_0_write_robId;
  assign integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid = Lsu2Plugin_setup_regfilePorts_0_write_valid;
  assign integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address = Lsu2Plugin_setup_regfilePorts_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_0_bypass_port_data = Lsu2Plugin_setup_regfilePorts_0_write_data;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_valid = (ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid != 1'b0);
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_address = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_data = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  assign integer_RegFilePlugin_logic_writeMerges_1_bus_robId = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId;
  assign integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid;
  assign integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_1_bypass_port_data = ALU0_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  assign integer_RegFilePlugin_logic_writeMerges_2_bus_valid = (ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_valid != 1'b0);
  assign integer_RegFilePlugin_logic_writeMerges_2_bus_address = ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_2_bus_data = ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  assign integer_RegFilePlugin_logic_writeMerges_2_bus_robId = ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_robId;
  assign integer_RegFilePlugin_logic_writeMerges_2_bypass_port_valid = ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_valid;
  assign integer_RegFilePlugin_logic_writeMerges_2_bypass_port_address = ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_2_bypass_port_data = ALU1_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  assign integer_RegFilePlugin_logic_writeMerges_3_bus_valid = (EU0_ExecutionUnitBase_pipeline_writeBack_0_write_valid != 1'b0);
  assign integer_RegFilePlugin_logic_writeMerges_3_bus_address = EU0_ExecutionUnitBase_pipeline_writeBack_0_write_address;
  assign integer_RegFilePlugin_logic_writeMerges_3_bus_data = EU0_ExecutionUnitBase_pipeline_writeBack_0_write_data;
  assign integer_RegFilePlugin_logic_writeMerges_3_bus_robId = EU0_ExecutionUnitBase_pipeline_writeBack_0_write_robId;
  assign EU0_ExecutionUnitBase_pipeline_writeBack_0_write_ready = 1'b1;
  always @(*) begin
    ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
    if(when_RegFilePlugin_l322) begin
      ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2;
    end
  end

  always @(*) begin
    ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
    if(when_RegFilePlugin_l322_1) begin
      ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2;
    end
  end

  always @(*) begin
    ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_2_data;
    if(when_RegFilePlugin_l322_2) begin
      ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2;
    end
  end

  always @(*) begin
    ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_3_data;
    if(when_RegFilePlugin_l322_3) begin
      ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2;
    end
  end

  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_4_data;
    if(when_RegFilePlugin_l322_4) begin
      EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_2;
    end
  end

  always @(*) begin
    EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_5_data;
    if(when_RegFilePlugin_l322_5) begin
      EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_2;
    end
  end

  assign _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1 = (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address));
  assign when_RegFilePlugin_l322 = ({_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1,{_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data,(integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address))}} != 3'b000);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address));
  assign _zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1 = (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address));
  assign when_RegFilePlugin_l322_1 = ({_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1,{_zz_ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data,(integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == ALU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address))}} != 3'b000);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address));
  assign _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1 = (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_address == ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address));
  assign when_RegFilePlugin_l322_2 = ({_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1,{_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data,(integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address))}} != 3'b000);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address));
  assign _zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1 = (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_address == ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address));
  assign when_RegFilePlugin_l322_3 = ({_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1,{_zz_ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data,(integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == ALU1_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address))}} != 3'b000);
  assign _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data = (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address));
  assign _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1 = (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address));
  assign when_RegFilePlugin_l322_4 = ({_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data_1,{_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_data,(integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS1_address))}} != 3'b000);
  assign _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data = (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_1_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address));
  assign _zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1 = (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_2_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address));
  assign when_RegFilePlugin_l322_5 = ({_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data_1,{_zz_EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_data,(integer_RegFilePlugin_logic_writeMerges_0_bypass_port_valid && (integer_RegFilePlugin_logic_writeMerges_0_bypass_port_address == EU0_ExecutionUnitBase_pipeline_rfReads_integer_RS2_address))}} != 3'b000);
  assign integer_write_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  assign integer_write_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  assign integer_write_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  assign integer_write_0_robId = integer_RegFilePlugin_logic_writeMerges_0_bus_robId;
  assign integer_write_1_valid = integer_RegFilePlugin_logic_writeMerges_1_bus_valid;
  assign integer_write_1_address = integer_RegFilePlugin_logic_writeMerges_1_bus_address;
  assign integer_write_1_data = integer_RegFilePlugin_logic_writeMerges_1_bus_data;
  assign integer_write_1_robId = integer_RegFilePlugin_logic_writeMerges_1_bus_robId;
  assign integer_write_2_valid = integer_RegFilePlugin_logic_writeMerges_2_bus_valid;
  assign integer_write_2_address = integer_RegFilePlugin_logic_writeMerges_2_bus_address;
  assign integer_write_2_data = integer_RegFilePlugin_logic_writeMerges_2_bus_data;
  assign integer_write_2_robId = integer_RegFilePlugin_logic_writeMerges_2_bus_robId;
  assign integer_write_3_valid = integer_RegFilePlugin_logic_writeMerges_3_bus_valid;
  assign integer_write_3_address = integer_RegFilePlugin_logic_writeMerges_3_bus_address;
  assign integer_write_3_data = integer_RegFilePlugin_logic_writeMerges_3_bus_data;
  assign integer_write_3_robId = integer_RegFilePlugin_logic_writeMerges_3_bus_robId;
  assign AguPlugin_setup_port_payload_earlySample = EU0_ExecutionUnitBase_pipeline_fetch_0_ready;
  assign AguPlugin_setup_port_payload_earlyPc = EU0_ExecutionUnitBase_pipeline_fetch_0_PC;
  assign RobPlugin_logic_completionMem_targetWrite_valid = FrontendPlugin_allocated_isFireing;
  assign RobPlugin_logic_completionMem_targetWrite_payload_address = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign RobPlugin_logic_completionMem_init_0_robId = {_zz_RobPlugin_logic_completionMem_init_0_robId,1'b0};
  always @(*) begin
    RobPlugin_logic_completionMem_targetWrite_payload_data[0] = ((((((_zz_RobPlugin_logic_completionMem_hits_0_port0[0] ^ _zz_RobPlugin_logic_completionMem_hits_1_port0[0]) ^ _zz_RobPlugin_logic_completionMem_hits_2_port0[0]) ^ _zz_RobPlugin_logic_completionMem_hits_3_port0[0]) ^ _zz_RobPlugin_logic_completionMem_hits_4_port0[0]) ^ _zz_RobPlugin_logic_completionMem_hits_5_port0[0]) ^ _zz_RobPlugin_logic_completionMem_hits_6_port0[0]);
    RobPlugin_logic_completionMem_targetWrite_payload_data[1] = ((((((_zz_RobPlugin_logic_completionMem_hits_0_port1[0] ^ _zz_RobPlugin_logic_completionMem_hits_1_port1[0]) ^ _zz_RobPlugin_logic_completionMem_hits_2_port1[0]) ^ _zz_RobPlugin_logic_completionMem_hits_3_port1[0]) ^ _zz_RobPlugin_logic_completionMem_hits_4_port1[0]) ^ _zz_RobPlugin_logic_completionMem_hits_5_port1[0]) ^ _zz_RobPlugin_logic_completionMem_hits_6_port1[0]);
  end

  assign RobPlugin_logic_completionMem_init_1_robId = {_zz_RobPlugin_logic_completionMem_init_1_robId,1'b1};
  assign RobPlugin_logic_completionMem_reads_0_targetRead_data = _zz_RobPlugin_logic_completionMem_target_port1;
  assign RobPlugin_logic_completionMem_reads_0_targetRead_address = (CommitPlugin_setup_robLineMask_line >>> 1'd1);
  assign _zz_CommitPlugin_setup_robLineMask_mask = {_zz__zz_CommitPlugin_setup_robLineMask_mask,1'b0};
  always @(*) begin
    CommitPlugin_setup_robLineMask_mask[0] = (((((((_zz_RobPlugin_logic_completionMem_hits_0_port4[0] ^ _zz_RobPlugin_logic_completionMem_hits_1_port4[0]) ^ _zz_RobPlugin_logic_completionMem_hits_2_port4[0]) ^ _zz_RobPlugin_logic_completionMem_hits_3_port4[0]) ^ _zz_RobPlugin_logic_completionMem_hits_4_port4[0]) ^ _zz_RobPlugin_logic_completionMem_hits_5_port4[0]) ^ _zz_RobPlugin_logic_completionMem_hits_6_port4[0]) != RobPlugin_logic_completionMem_reads_0_targetRead_data[0]);
    CommitPlugin_setup_robLineMask_mask[1] = (((((((_zz_RobPlugin_logic_completionMem_hits_0_port5[0] ^ _zz_RobPlugin_logic_completionMem_hits_1_port5[0]) ^ _zz_RobPlugin_logic_completionMem_hits_2_port5[0]) ^ _zz_RobPlugin_logic_completionMem_hits_3_port5[0]) ^ _zz_RobPlugin_logic_completionMem_hits_4_port5[0]) ^ _zz_RobPlugin_logic_completionMem_hits_5_port5[0]) ^ _zz_RobPlugin_logic_completionMem_hits_6_port5[0]) != RobPlugin_logic_completionMem_reads_0_targetRead_data[1]);
    if(when_RobPlugin_l118) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_1) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_2) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_3) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_4) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_5) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_6) begin
      CommitPlugin_setup_robLineMask_mask[0] = 1'b1;
    end
    if(when_RobPlugin_l118_7) begin
      CommitPlugin_setup_robLineMask_mask[1] = 1'b1;
    end
    if(when_RobPlugin_l118_8) begin
      CommitPlugin_setup_robLineMask_mask[1] = 1'b1;
    end
    if(when_RobPlugin_l118_9) begin
      CommitPlugin_setup_robLineMask_mask[1] = 1'b1;
    end
    if(when_RobPlugin_l118_10) begin
      CommitPlugin_setup_robLineMask_mask[1] = 1'b1;
    end
    if(when_RobPlugin_l118_11) begin
      CommitPlugin_setup_robLineMask_mask[1] = 1'b1;
    end
    if(when_RobPlugin_l118_12) begin
      CommitPlugin_setup_robLineMask_mask[1] = 1'b1;
    end
    if(when_RobPlugin_l118_13) begin
      CommitPlugin_setup_robLineMask_mask[1] = 1'b1;
    end
    if(when_RobPlugin_l123) begin
      CommitPlugin_setup_robLineMask_mask = 2'b00;
    end
  end

  assign _zz_CommitPlugin_setup_robLineMask_mask_1 = {_zz__zz_CommitPlugin_setup_robLineMask_mask_1,1'b1};
  assign _zz_when_RobPlugin_l118 = {_zz__zz_when_RobPlugin_l118,1'b0};
  assign when_RobPlugin_l118 = (Lsu2Plugin_setup_sharedCompletion_valid && (Lsu2Plugin_setup_sharedCompletion_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l118_1 = (Lsu2Plugin_setup_specialCompletion_valid && (Lsu2Plugin_setup_specialCompletion_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l118_2 = (ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid && (ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l118_3 = (ALU0_ExecutionUnitBase_pipeline_completion_1_port_valid && (ALU0_ExecutionUnitBase_pipeline_completion_1_port_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l118_4 = (ALU1_ExecutionUnitBase_pipeline_completion_0_port_valid && (ALU1_ExecutionUnitBase_pipeline_completion_0_port_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l118_5 = (ALU1_ExecutionUnitBase_pipeline_completion_1_port_valid && (ALU1_ExecutionUnitBase_pipeline_completion_1_port_payload_id == _zz_when_RobPlugin_l118));
  assign when_RobPlugin_l118_6 = (EU0_ExecutionUnitBase_pipeline_completion_0_port_valid && (EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id == _zz_when_RobPlugin_l118));
  assign _zz_when_RobPlugin_l118_1 = {_zz__zz_when_RobPlugin_l118_1,1'b1};
  assign when_RobPlugin_l118_7 = (Lsu2Plugin_setup_sharedCompletion_valid && (Lsu2Plugin_setup_sharedCompletion_payload_id == _zz_when_RobPlugin_l118_1));
  assign when_RobPlugin_l118_8 = (Lsu2Plugin_setup_specialCompletion_valid && (Lsu2Plugin_setup_specialCompletion_payload_id == _zz_when_RobPlugin_l118_1));
  assign when_RobPlugin_l118_9 = (ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid && (ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id == _zz_when_RobPlugin_l118_1));
  assign when_RobPlugin_l118_10 = (ALU0_ExecutionUnitBase_pipeline_completion_1_port_valid && (ALU0_ExecutionUnitBase_pipeline_completion_1_port_payload_id == _zz_when_RobPlugin_l118_1));
  assign when_RobPlugin_l118_11 = (ALU1_ExecutionUnitBase_pipeline_completion_0_port_valid && (ALU1_ExecutionUnitBase_pipeline_completion_0_port_payload_id == _zz_when_RobPlugin_l118_1));
  assign when_RobPlugin_l118_12 = (ALU1_ExecutionUnitBase_pipeline_completion_1_port_valid && (ALU1_ExecutionUnitBase_pipeline_completion_1_port_payload_id == _zz_when_RobPlugin_l118_1));
  assign when_RobPlugin_l118_13 = (EU0_ExecutionUnitBase_pipeline_completion_0_port_valid && (EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id == _zz_when_RobPlugin_l118_1));
  assign when_RobPlugin_l123 = (FrontendPlugin_allocated_isFireing && (FrontendPlugin_allocated_ROB_ID == CommitPlugin_setup_robLineMask_line));
  assign _zz_CommitPlugin_logic_commit_active = (CommitPlugin_logic_ptr_commit[5 : 0] >>> 1'd1);
  assign _zz_CommitPlugin_logic_commit_active_1 = _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port1;
  assign _zz_CommitPlugin_logic_commit_active_2 = _zz__zz_CommitPlugin_logic_commit_active_2[1 : 0];
  assign _zz_integer_RfAllocationPlugin_logic_push_mask_0 = (CommitPlugin_logic_free_port_payload_robId >>> 1'd1);
  assign _zz_integer_RfAllocationPlugin_logic_push_mask_0_1 = _zz_RobPlugin_logic_storage_Frontend_DISPATCH_MASK_banks_0_port2;
  assign _zz_integer_RfAllocationPlugin_logic_push_mask_0_2 = _zz__zz_integer_RfAllocationPlugin_logic_push_mask_0_2[1 : 0];
  assign integer_RfAllocationPlugin_logic_push_mask_0 = _zz_integer_RfAllocationPlugin_logic_push_mask_0_2[0];
  assign integer_RfAllocationPlugin_logic_push_mask_1 = _zz_integer_RfAllocationPlugin_logic_push_mask_0_2[1];
  assign _zz_224 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_commit_pc_0 = (CommitPlugin_logic_commit_event_robId >>> 1'd1);
  assign _zz_commit_pc_0_1 = _zz__zz_commit_pc_0_1[63 : 0];
  assign _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc = (CommitPlugin_logic_commit_reschedulePort_payload_robId >>> 1'd1);
  assign _zz_PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc_1 = {_zz_RobPlugin_logic_storage_PC_banks_1_port2[31 : 0],_zz_RobPlugin_logic_storage_PC_banks_0_port2[31 : 0]};
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PC = (ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PC = (ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC = (EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_PC_1 = {_zz_RobPlugin_logic_storage_PC_banks_1_port4[31 : 0],_zz_RobPlugin_logic_storage_PC_banks_0_port4[31 : 0]};
  assign _zz_235 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0 = (CommitPlugin_logic_commit_event_robId >>> 1'd1);
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1 = _zz__zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1[1 : 0];
  assign integer_RfTranslationPlugin_logic_onCommit_writeRd_0 = _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1[0];
  assign integer_RfTranslationPlugin_logic_onCommit_writeRd_1 = _zz_integer_RfTranslationPlugin_logic_onCommit_writeRd_0_1[1];
  assign _zz_integer_RfAllocationPlugin_logic_push_writeRd_0 = (CommitPlugin_logic_free_port_payload_robId >>> 1'd1);
  assign _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1 = _zz__zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1[1 : 0];
  assign integer_RfAllocationPlugin_logic_push_writeRd_0 = _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1[0];
  assign integer_RfAllocationPlugin_logic_push_writeRd_1 = _zz_integer_RfAllocationPlugin_logic_push_writeRd_0_1[1];
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = (ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = (ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD = (EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD_1 = {_zz_RobPlugin_logic_storage_WRITE_RD_banks_1_port4[0],_zz_RobPlugin_logic_storage_WRITE_RD_banks_0_port4[0]};
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0 = (CommitPlugin_logic_commit_event_robId >>> 1'd1);
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_1 = _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port1;
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2 = _zz__zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2[11 : 0];
  assign integer_RfTranslationPlugin_logic_onCommit_physRd_0 = _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2[5 : 0];
  assign integer_RfTranslationPlugin_logic_onCommit_physRd_1 = _zz_integer_RfTranslationPlugin_logic_onCommit_physRd_0_2[11 : 6];
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0 = (CommitPlugin_logic_free_port_payload_robId >>> 1'd1);
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_1 = _zz_RobPlugin_logic_storage_PHYS_RD_banks_0_port2;
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2 = _zz__zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2[11 : 0];
  assign integer_RfAllocationPlugin_logic_push_physicalRdNew_0 = _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2[5 : 0];
  assign integer_RfAllocationPlugin_logic_push_physicalRdNew_1 = _zz_integer_RfAllocationPlugin_logic_push_physicalRdNew_0_2[11 : 6];
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0 = (CommitPlugin_logic_commit_event_robId >>> 1'd1);
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_1 = _zz_RobPlugin_logic_storage_ARCH_RD_banks_0_port1;
  assign _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2 = _zz__zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2[9 : 0];
  assign integer_RfTranslationPlugin_logic_onCommit_archRd_0 = _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2[4 : 0];
  assign integer_RfTranslationPlugin_logic_onCommit_archRd_1 = _zz_integer_RfTranslationPlugin_logic_onCommit_archRd_0_2[9 : 5];
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0 = (CommitPlugin_logic_free_port_payload_robId >>> 1'd1);
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_1 = _zz_RobPlugin_logic_storage_PHYS_RD_FREE_banks_0_port1;
  assign _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2 = _zz__zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2[11 : 0];
  assign integer_RfAllocationPlugin_logic_push_physicalRdOld_0 = _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2[5 : 0];
  assign integer_RfAllocationPlugin_logic_push_physicalRdOld_1 = _zz_integer_RfAllocationPlugin_logic_push_physicalRdOld_0_2[11 : 6];
  assign _zz_BranchContextPlugin_logic_onCommit_isBranch_0 = (CommitPlugin_logic_commit_event_robId >>> 1'd1);
  assign _zz_BranchContextPlugin_logic_onCommit_isBranch_0_1 = _zz_RobPlugin_logic_storage_BRANCH_SEL_banks_0_port1;
  assign _zz_BranchContextPlugin_logic_onCommit_isBranch_0_2 = _zz__zz_BranchContextPlugin_logic_onCommit_isBranch_0_2[1 : 0];
  assign BranchContextPlugin_logic_onCommit_isBranch_0 = _zz_BranchContextPlugin_logic_onCommit_isBranch_0_2[0];
  assign BranchContextPlugin_logic_onCommit_isBranch_1 = _zz_BranchContextPlugin_logic_onCommit_isBranch_0_2[1];
  assign _zz_255 = (FrontendPlugin_dispatch_ROB_ID >>> 1'd1);
  assign _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0 = (CommitPlugin_logic_commit_event_robId >>> 1'd1);
  assign _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1 = _zz__zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1[1 : 0];
  assign HistoryPlugin_logic_onCommit_isConditionalBranch_0 = _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1[0];
  assign HistoryPlugin_logic_onCommit_isConditionalBranch_1 = _zz_HistoryPlugin_logic_onCommit_isConditionalBranch_0_1[1];
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch = (CommitPlugin_logic_reschedule_reschedulePort_payload_robId >>> 1'd1);
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_isConditionalBranch_1 = {_zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_1_port2[0],_zz_RobPlugin_logic_storage_Prediction_IS_BRANCH_banks_0_port2[0]};
  assign _zz_io_read_0_cmd_payload = (CommitPlugin_logic_commit_event_robId >>> 1'd1);
  assign _zz_HistoryPlugin_logic_onCommit_isTaken_0 = {RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_1_rsp[0],RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_0_rsp[0]};
  assign HistoryPlugin_logic_onCommit_isTaken_0 = _zz_HistoryPlugin_logic_onCommit_isTaken_0[0];
  assign HistoryPlugin_logic_onCommit_isTaken_1 = _zz_HistoryPlugin_logic_onCommit_isTaken_0[1];
  assign _zz_262 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory = (CommitPlugin_logic_reschedule_reschedulePort_payload_robId >>> 1'd1);
  assign _zz_HistoryPlugin_logic_update_rescheduleFlush_instHistory_1 = {_zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_1_port1[23 : 0],_zz_RobPlugin_logic_storage_BRANCH_HISTORY_banks_0_port1[23 : 0]};
  assign _zz_267 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_DecoderPredictionPlugin_logic_ras_healPush = (CommitPlugin_logic_reschedule_reschedulePort_payload_robId >>> 1'd1);
  assign _zz_DecoderPredictionPlugin_logic_ras_healPush_1 = {_zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_1_port1[3 : 0],_zz_RobPlugin_logic_storage_DecoderPredictionPlugin_RAS_PUSH_PTR_banks_0_port1[3 : 0]};
  assign _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0 = (CommitPlugin_logic_commit_event_robId >>> 1'd1);
  assign _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_1 = _zz_RobPlugin_logic_storage_LQ_ALLOC_banks_0_port1;
  assign _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2 = _zz__zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2[1 : 0];
  assign Lsu2Plugin_logic_lq_onCommit_lqAlloc_0 = _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2[0];
  assign Lsu2Plugin_logic_lq_onCommit_lqAlloc_1 = _zz_Lsu2Plugin_logic_lq_onCommit_lqAlloc_0_2[1];
  assign _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0 = (CommitPlugin_logic_commit_event_robId >>> 1'd1);
  assign _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_1 = _zz_RobPlugin_logic_storage_SQ_ALLOC_banks_0_port1;
  assign _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2 = _zz__zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2[1 : 0];
  assign Lsu2Plugin_logic_sq_onCommit_sqAlloc_0 = _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2[0];
  assign Lsu2Plugin_logic_sq_onCommit_sqAlloc_1 = _zz_Lsu2Plugin_logic_sq_onCommit_sqAlloc_0_2[1];
  assign _zz_276 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = (ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = (ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP = (EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP_1 = {_zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_1_port2[31 : 0],_zz_RobPlugin_logic_storage_Frontend_MICRO_OP_banks_0_port2[31 : 0]};
  assign _zz_283 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0 = (ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_0 = (ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_288 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = (ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = (ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0 = (EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_0_1 = {_zz_RobPlugin_logic_storage_READ_RS_0_banks_1_port2[0],_zz_RobPlugin_logic_storage_READ_RS_0_banks_0_port2[0]};
  assign _zz_295 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1 = (ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RS_1 = (ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_300 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = (ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = (ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1 = (EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_READ_RS_1_1 = {_zz_RobPlugin_logic_storage_READ_RS_1_banks_1_port2[0],_zz_RobPlugin_logic_storage_READ_RS_1_banks_0_port2[0]};
  assign _zz_307 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID = (ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID = (ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_312 = (FrontendPlugin_dispatch_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID = (EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID_1 = {_zz_RobPlugin_logic_storage_LSU_ID_banks_1_port1[4 : 0],_zz_RobPlugin_logic_storage_LSU_ID_banks_0_port1[4 : 0]};
  assign _zz_317 = (FrontendPlugin_allocated_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB = (EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID >>> 1'd1);
  assign _zz_EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB_1 = {_zz_RobPlugin_logic_storage_ROB_MSB_banks_1_port1[0 : 0],_zz_RobPlugin_logic_storage_ROB_MSB_banks_0_port1[0 : 0]};
  assign RobPlugin_logic_whitebox_completionsPorts_0_valid = Lsu2Plugin_setup_sharedCompletion_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_0_payload_id = Lsu2Plugin_setup_sharedCompletion_payload_id;
  assign RobPlugin_logic_whitebox_completionsPorts_1_valid = Lsu2Plugin_setup_specialCompletion_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_1_payload_id = Lsu2Plugin_setup_specialCompletion_payload_id;
  assign RobPlugin_logic_whitebox_completionsPorts_2_valid = ALU0_ExecutionUnitBase_pipeline_completion_0_port_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_2_payload_id = ALU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  assign RobPlugin_logic_whitebox_completionsPorts_3_valid = ALU0_ExecutionUnitBase_pipeline_completion_1_port_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_3_payload_id = ALU0_ExecutionUnitBase_pipeline_completion_1_port_payload_id;
  assign RobPlugin_logic_whitebox_completionsPorts_4_valid = ALU1_ExecutionUnitBase_pipeline_completion_0_port_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_4_payload_id = ALU1_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  assign RobPlugin_logic_whitebox_completionsPorts_5_valid = ALU1_ExecutionUnitBase_pipeline_completion_1_port_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_5_payload_id = ALU1_ExecutionUnitBase_pipeline_completion_1_port_payload_id;
  assign RobPlugin_logic_whitebox_completionsPorts_6_valid = EU0_ExecutionUnitBase_pipeline_completion_0_port_valid;
  assign RobPlugin_logic_whitebox_completionsPorts_6_payload_id = EU0_ExecutionUnitBase_pipeline_completion_0_port_payload_id;
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_valid = (((FrontendPlugin_dispatch_isFireing && FrontendPlugin_dispatch_WRITE_RD_0) && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_writes_0_payload_robId = (FrontendPlugin_dispatch_ROB_ID | 6'h00);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_writes_1_valid = (((FrontendPlugin_dispatch_isFireing && FrontendPlugin_dispatch_WRITE_RD_1) && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1) && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_writes_1_payload_robId = (FrontendPlugin_dispatch_ROB_ID | 6'h01);
  always @(*) begin
    RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_valid = (DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid && 1'b1);
    if(RfDependencyPlugin_logic_forRf_integer_init_busy) begin
      RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_valid = 1'b1;
    end
  end

  always @(*) begin
    RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_payload_physical = DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical;
    if(RfDependencyPlugin_logic_forRf_integer_init_busy) begin
      RfDependencyPlugin_logic_forRf_integer_impl_io_commits_0_payload_physical = RfDependencyPlugin_logic_forRf_integer_init_counter[5:0];
    end
  end

  assign RfDependencyPlugin_logic_forRf_integer_impl_io_commits_1_valid = (DispatchPlugin_logic_pop_1_wake_L0_bypassed_valid && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_commits_2_valid = (Lsu2Plugin_logic_sharedPip_hitSpeculation_wakeRf_valid && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_commits_3_valid = (Lsu2Plugin_logic_sharedPip_ctrl_wakeRf_valid && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_commits_4_valid = (Lsu2Plugin_logic_special_wakeRf_valid && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_commits_5_valid = (EU0_ExecutionUnitBase_pipeline_wakeRf_logic_0_rf_valid && 1'b1);
  assign RfDependencyPlugin_logic_forRf_integer_init_busy = (! RfDependencyPlugin_logic_forRf_integer_init_counter[6]);
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_cmd_valid = ((FrontendPlugin_dispatch_valid && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && FrontendPlugin_dispatch_READ_RS_0_0);
  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = 1'bx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_enable;
  end

  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0 = 6'bxxxxxx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_0_rsp_payload_rob;
  end

  always @(*) begin
    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0;
    if(when_RfDependencyPlugin_l241) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = 1'b0;
    end
    if(when_RfDependencyPlugin_l241_1) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = 1'b0;
    end
    if(when_RfDependencyPlugin_l245) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 = 1'b0;
    end
  end

  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_0;
  assign when_RfDependencyPlugin_l241 = ((DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_0_0)) && 1'b1);
  assign when_RfDependencyPlugin_l241_1 = ((DispatchPlugin_logic_pop_1_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_1_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_0_0)) && 1'b1);
  assign when_RfDependencyPlugin_l245 = (! FrontendPlugin_dispatch_READ_RS_0_0);
  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_0 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_0 && (! FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_0_0));
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_cmd_valid = ((FrontendPlugin_dispatch_valid && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && FrontendPlugin_dispatch_READ_RS_1_0);
  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = 1'bx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_enable;
  end

  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0 = 6'bxxxxxx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_1_rsp_payload_rob;
  end

  always @(*) begin
    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0;
    if(when_RfDependencyPlugin_l241_2) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = 1'b0;
    end
    if(when_RfDependencyPlugin_l241_3) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = 1'b0;
    end
    if(when_RfDependencyPlugin_l245_1) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 = 1'b0;
    end
  end

  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_0;
  assign when_RfDependencyPlugin_l241_2 = ((DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_1_0)) && 1'b1);
  assign when_RfDependencyPlugin_l241_3 = ((DispatchPlugin_logic_pop_1_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_1_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_1_0)) && 1'b1);
  assign when_RfDependencyPlugin_l245_1 = (! FrontendPlugin_dispatch_READ_RS_1_0);
  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_0 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_0 && (! FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_1_0));
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_cmd_valid = ((FrontendPlugin_dispatch_valid && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1) && FrontendPlugin_dispatch_READ_RS_0_1);
  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1 = 1'bx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_rsp_payload_enable;
  end

  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_1 = 6'bxxxxxx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_1 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_2_rsp_payload_rob;
  end

  always @(*) begin
    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1;
    if(when_RfDependencyPlugin_l235) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1 = 1'b1;
    end
    if(when_RfDependencyPlugin_l241_4) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1 = 1'b0;
    end
    if(when_RfDependencyPlugin_l241_5) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1 = 1'b0;
    end
    if(when_RfDependencyPlugin_l245_2) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1 = 1'b0;
    end
  end

  always @(*) begin
    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_1 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_1;
    if(when_RfDependencyPlugin_l235) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ID_1 = (FrontendPlugin_dispatch_ROB_ID | 6'h00);
    end
  end

  assign when_RfDependencyPlugin_l235 = (((FrontendPlugin_dispatch_WRITE_RD_0 && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && 1'b1) && (FrontendPlugin_dispatch_ARCH_RD_0 == FrontendPlugin_dispatch_ARCH_RS_0_1));
  assign when_RfDependencyPlugin_l241_4 = ((DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_0_1)) && 1'b1);
  assign when_RfDependencyPlugin_l241_5 = ((DispatchPlugin_logic_pop_1_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_1_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_0_1)) && 1'b1);
  assign when_RfDependencyPlugin_l245_2 = (! FrontendPlugin_dispatch_READ_RS_0_1);
  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_1 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_0_ENABLE_UNSKIPED_1 && (! FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_0_1));
  assign RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_cmd_valid = ((FrontendPlugin_dispatch_valid && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1) && FrontendPlugin_dispatch_READ_RS_1_1);
  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1 = 1'bx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_rsp_payload_enable;
  end

  always @(*) begin
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_1 = 6'bxxxxxx;
    _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_1 = RfDependencyPlugin_logic_forRf_integer_impl_io_reads_3_rsp_payload_rob;
  end

  always @(*) begin
    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1;
    if(when_RfDependencyPlugin_l235_1) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1 = 1'b1;
    end
    if(when_RfDependencyPlugin_l241_6) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1 = 1'b0;
    end
    if(when_RfDependencyPlugin_l241_7) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1 = 1'b0;
    end
    if(when_RfDependencyPlugin_l245_3) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1 = 1'b0;
    end
  end

  always @(*) begin
    FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_1 = _zz_FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_1;
    if(when_RfDependencyPlugin_l235_1) begin
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ID_1 = (FrontendPlugin_dispatch_ROB_ID | 6'h00);
    end
  end

  assign when_RfDependencyPlugin_l235_1 = (((FrontendPlugin_dispatch_WRITE_RD_0 && FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0) && 1'b1) && (FrontendPlugin_dispatch_ARCH_RD_0 == FrontendPlugin_dispatch_ARCH_RS_1_1));
  assign when_RfDependencyPlugin_l241_6 = ((DispatchPlugin_logic_pop_0_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_0_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_1_1)) && 1'b1);
  assign when_RfDependencyPlugin_l241_7 = ((DispatchPlugin_logic_pop_1_wake_L0_bypassed_valid && (DispatchPlugin_logic_pop_1_wake_L0_bypassed_payload_physical == FrontendPlugin_dispatch_PHYS_RS_1_1)) && 1'b1);
  assign when_RfDependencyPlugin_l245_3 = (! FrontendPlugin_dispatch_READ_RS_1_1);
  assign FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_1 = (FrontendPlugin_dispatch_RfDependencyPlugin_setup_waits_1_ENABLE_UNSKIPED_1 && (! FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_1_1));
  assign FrontendPlugin_isBusy = ({FrontendPlugin_dispatch_valid,{FrontendPlugin_allocated_valid,{FrontendPlugin_serialized_valid,{FrontendPlugin_decoded_valid,FrontendPlugin_decompressed_valid}}}} != 5'h00);
  assign FrontendPlugin_isBusyAfterDecode = ({FrontendPlugin_dispatch_valid,{FrontendPlugin_allocated_valid,FrontendPlugin_serialized_valid}} != 3'b000);
  assign FrontendPlugin_dispatch_isFlushed = CommitPlugin_logic_reschedule_reschedulePort_valid;
  assign FrontendPlugin_allocated_isFlushed = CommitPlugin_logic_reschedule_reschedulePort_valid;
  assign when_Connection_l66 = ({CommitPlugin_logic_reschedule_reschedulePort_valid,(DecoderPredictionPlugin_setup_decodeJump_valid && FrontendPlugin_serialized_ready)} != 2'b00);
  assign FrontendPlugin_serialized_isFlushed = when_Connection_l66;
  assign _zz_FrontendPlugin_decompressed_isFlushed = ({when_Connection_l66,_zz_FrontendPlugin_decoded_isFlushingRoot} != 2'b00);
  assign FrontendPlugin_decoded_isFlushed = _zz_FrontendPlugin_decompressed_isFlushed;
  assign FrontendPlugin_decompressed_isFlushed = _zz_FrontendPlugin_decompressed_isFlushed;
  assign FrontendPlugin_aligned_isFlushed = _zz_FrontendPlugin_decompressed_isFlushed;
  assign FrontendPlugin_decoded_isFlushingRoot = (_zz_FrontendPlugin_decoded_isFlushingRoot != 1'b0);
  assign FrontendPlugin_dispatch_isFlushingRoot = (CommitPlugin_logic_reschedule_reschedulePort_valid != 1'b0);
  assign FrontendPlugin_serialized_isForked = (_zz_FrontendPlugin_serialized_isForked && FrontendPlugin_serialized_ready_output);
  assign FrontendPlugin_aligned_ready = FrontendPlugin_aligned_ready_output;
  assign FrontendPlugin_decompressed_ready = FrontendPlugin_decompressed_ready_output;
  always @(*) begin
    _zz_FrontendPlugin_serialized_valid = FrontendPlugin_decoded_valid;
    if(FrontendPlugin_decoded_isFlushingRoot) begin
      _zz_FrontendPlugin_serialized_valid = 1'b0;
    end
    if(when_Pipeline_l278_6) begin
      _zz_FrontendPlugin_serialized_valid = 1'b0;
    end
  end

  always @(*) begin
    FrontendPlugin_decoded_ready = FrontendPlugin_decoded_ready_output;
    if(when_Pipeline_l278_6) begin
      FrontendPlugin_decoded_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_6 = ({FrontendPlugin_decoded_haltRequest_DecoderPlugin_l323,FrontendPlugin_decoded_haltRequest_DecoderPlugin_l322} != 2'b00);
  assign _zz_FrontendPlugin_serialized_isForked = FrontendPlugin_serialized_valid;
  always @(*) begin
    FrontendPlugin_serialized_ready = FrontendPlugin_serialized_ready_output;
    if(when_Pipeline_l285) begin
      FrontendPlugin_serialized_ready = 1'b0;
    end
  end

  assign when_Pipeline_l285 = (FrontendPlugin_serialized_forkRequest_DispatchPlugin_l90 != 1'b0);
  always @(*) begin
    _zz_FrontendPlugin_dispatch_valid = FrontendPlugin_allocated_valid;
    if(when_Pipeline_l278_7) begin
      _zz_FrontendPlugin_dispatch_valid = 1'b0;
    end
  end

  always @(*) begin
    FrontendPlugin_allocated_ready = FrontendPlugin_allocated_ready_output;
    if(when_Pipeline_l278_7) begin
      FrontendPlugin_allocated_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_7 = ({FrontendPlugin_allocated_haltRequest_FrontendPlugin_l67,{FrontendPlugin_allocated_haltRequest_CommitPlugin_l95,{FrontendPlugin_allocated_haltRequest_BranchContextPlugin_l107,FrontendPlugin_allocated_haltRequest_RfAllocationPlugin_l55}}} != 4'b0000);
  always @(*) begin
    FrontendPlugin_dispatch_ready = 1'b1;
    if(when_Pipeline_l278_8) begin
      FrontendPlugin_dispatch_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_8 = ({FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l196,{FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l195,{FrontendPlugin_dispatch_haltRequest_DispatchPlugin_l187,{FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l1834,FrontendPlugin_dispatch_haltRequest_Lsu2Plugin_l620}}}} != 5'h00);
  assign FrontendPlugin_serialized_ready_output = FrontendPlugin_allocated_ready;
  assign FrontendPlugin_allocated_valid = _zz_FrontendPlugin_serialized_isForked;
  assign FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0 = FrontendPlugin_serialized_Frontend_DISPATCH_MASK_0_overloaded;
  assign FrontendPlugin_allocated_Frontend_DISPATCH_MASK_1 = FrontendPlugin_serialized_Frontend_DISPATCH_MASK_1_overloaded;
  assign FrontendPlugin_allocated_DispatchPlugin_FENCE_OLDER_0 = FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_0;
  assign FrontendPlugin_allocated_Frontend_MICRO_OP_0 = FrontendPlugin_serialized_Frontend_MICRO_OP_0;
  assign FrontendPlugin_allocated_DispatchPlugin_FENCE_YOUNGER_0 = FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_0;
  assign FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_0_0 = FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_0;
  assign FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_1_0 = FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_0;
  assign FrontendPlugin_allocated_DispatchPlugin_FENCE_OLDER_1 = FrontendPlugin_serialized_DispatchPlugin_FENCE_OLDER_1;
  assign FrontendPlugin_allocated_Frontend_MICRO_OP_1 = FrontendPlugin_serialized_Frontend_MICRO_OP_1;
  assign FrontendPlugin_allocated_DispatchPlugin_FENCE_YOUNGER_1 = FrontendPlugin_serialized_DispatchPlugin_FENCE_YOUNGER_1;
  assign FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_0_1 = FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_0_1;
  assign FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_1_1 = FrontendPlugin_serialized_RfDependencyPlugin_setup_SKIP_1_1;
  assign FrontendPlugin_allocated_BRANCH_SEL_0 = FrontendPlugin_serialized_BRANCH_SEL_0;
  assign FrontendPlugin_allocated_BRANCH_EARLY_0_taken = FrontendPlugin_serialized_BRANCH_EARLY_0_taken;
  assign FrontendPlugin_allocated_BRANCH_EARLY_0_pc = FrontendPlugin_serialized_BRANCH_EARLY_0_pc;
  assign FrontendPlugin_allocated_DecoderPredictionPlugin_RAS_PUSH_PTR_0 = FrontendPlugin_serialized_DecoderPredictionPlugin_RAS_PUSH_PTR_0;
  assign FrontendPlugin_allocated_BRANCH_SEL_1 = FrontendPlugin_serialized_BRANCH_SEL_1;
  assign FrontendPlugin_allocated_BRANCH_EARLY_1_taken = FrontendPlugin_serialized_BRANCH_EARLY_1_taken;
  assign FrontendPlugin_allocated_BRANCH_EARLY_1_pc = FrontendPlugin_serialized_BRANCH_EARLY_1_pc;
  assign FrontendPlugin_allocated_DecoderPredictionPlugin_RAS_PUSH_PTR_1 = FrontendPlugin_serialized_DecoderPredictionPlugin_RAS_PUSH_PTR_1;
  assign FrontendPlugin_allocated_Prediction_IS_BRANCH_0 = FrontendPlugin_serialized_Prediction_IS_BRANCH_0;
  assign FrontendPlugin_allocated_Prediction_IS_BRANCH_1 = FrontendPlugin_serialized_Prediction_IS_BRANCH_1;
  assign FrontendPlugin_allocated_FETCH_ID_0 = FrontendPlugin_serialized_FETCH_ID_0;
  assign FrontendPlugin_allocated_FETCH_ID_1 = FrontendPlugin_serialized_FETCH_ID_1;
  assign FrontendPlugin_allocated_WRITE_RD_0 = FrontendPlugin_serialized_WRITE_RD_0;
  assign FrontendPlugin_allocated_WRITE_RD_1 = FrontendPlugin_serialized_WRITE_RD_1;
  assign FrontendPlugin_allocated_PC_0 = FrontendPlugin_serialized_PC_0;
  assign FrontendPlugin_allocated_PC_1 = FrontendPlugin_serialized_PC_1;
  assign FrontendPlugin_allocated_ARCH_RD_0 = FrontendPlugin_serialized_ARCH_RD_0;
  assign FrontendPlugin_allocated_ARCH_RD_1 = FrontendPlugin_serialized_ARCH_RD_1;
  assign FrontendPlugin_allocated_ARCH_RS_0_0 = FrontendPlugin_serialized_ARCH_RS_0_0;
  assign FrontendPlugin_allocated_READ_RS_0_0 = FrontendPlugin_serialized_READ_RS_0_0;
  assign FrontendPlugin_allocated_ARCH_RS_1_0 = FrontendPlugin_serialized_ARCH_RS_1_0;
  assign FrontendPlugin_allocated_READ_RS_1_0 = FrontendPlugin_serialized_READ_RS_1_0;
  assign FrontendPlugin_allocated_ARCH_RS_0_1 = FrontendPlugin_serialized_ARCH_RS_0_1;
  assign FrontendPlugin_allocated_READ_RS_0_1 = FrontendPlugin_serialized_READ_RS_0_1;
  assign FrontendPlugin_allocated_ARCH_RS_1_1 = FrontendPlugin_serialized_ARCH_RS_1_1;
  assign FrontendPlugin_allocated_READ_RS_1_1 = FrontendPlugin_serialized_READ_RS_1_1;
  assign FrontendPlugin_allocated_BRANCH_HISTORY_0 = FrontendPlugin_serialized_BRANCH_HISTORY_0;
  assign FrontendPlugin_allocated_BRANCH_HISTORY_1 = FrontendPlugin_serialized_BRANCH_HISTORY_1;
  assign FrontendPlugin_allocated_OP_ID = FrontendPlugin_serialized_OP_ID;
  assign FrontendPlugin_allocated_LQ_ALLOC_0 = FrontendPlugin_serialized_LQ_ALLOC_0;
  assign FrontendPlugin_allocated_LQ_ALLOC_1 = FrontendPlugin_serialized_LQ_ALLOC_1;
  assign FrontendPlugin_allocated_SQ_ALLOC_0 = FrontendPlugin_serialized_SQ_ALLOC_0;
  assign FrontendPlugin_allocated_SQ_ALLOC_1 = FrontendPlugin_serialized_SQ_ALLOC_1;
  assign FrontendPlugin_allocated_GSHARE_COUNTER_0_0 = FrontendPlugin_serialized_GSHARE_COUNTER_0_0;
  assign FrontendPlugin_allocated_GSHARE_COUNTER_0_1 = FrontendPlugin_serialized_GSHARE_COUNTER_0_1;
  assign FrontendPlugin_allocated_GSHARE_COUNTER_1_0 = FrontendPlugin_serialized_GSHARE_COUNTER_1_0;
  assign FrontendPlugin_allocated_GSHARE_COUNTER_1_1 = FrontendPlugin_serialized_GSHARE_COUNTER_1_1;
  assign FrontendPlugin_allocated_ALU0_ALU1_SEL_0 = FrontendPlugin_serialized_ALU0_ALU1_SEL_0;
  assign FrontendPlugin_allocated_EU0_SEL_0 = FrontendPlugin_serialized_EU0_SEL_0;
  assign FrontendPlugin_allocated_ALU0_ALU1_SEL_1 = FrontendPlugin_serialized_ALU0_ALU1_SEL_1;
  assign FrontendPlugin_allocated_EU0_SEL_1 = FrontendPlugin_serialized_EU0_SEL_1;
  always @(*) begin
    FrontendPlugin_allocated_ready_output = FrontendPlugin_dispatch_ready;
    if(when_Connection_l74_5) begin
      FrontendPlugin_allocated_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_5 = (! FrontendPlugin_dispatch_valid);
  assign FrontendPlugin_aligned_ready_output = FrontendPlugin_decompressed_ready;
  assign FrontendPlugin_decompressed_valid = FrontendPlugin_aligned_valid;
  assign FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_0 = FrontendPlugin_aligned_Frontend_INSTRUCTION_ALIGNED_0;
  assign FrontendPlugin_decompressed_Frontend_MASK_ALIGNED_0 = FrontendPlugin_aligned_Frontend_MASK_ALIGNED_0;
  assign FrontendPlugin_decompressed_PC_0 = FrontendPlugin_aligned_PC_0;
  assign FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_VALID_0 = FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_0;
  assign FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_PC_NEXT_0 = FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  assign FrontendPlugin_decompressed_BRANCH_HISTORY_0 = FrontendPlugin_aligned_BRANCH_HISTORY_0;
  assign FrontendPlugin_decompressed_GSHARE_COUNTER_0_0 = FrontendPlugin_aligned_GSHARE_COUNTER_0_0;
  assign FrontendPlugin_decompressed_GSHARE_COUNTER_0_1 = FrontendPlugin_aligned_GSHARE_COUNTER_0_1;
  assign FrontendPlugin_decompressed_FETCH_ID_0 = FrontendPlugin_aligned_FETCH_ID_0;
  assign FrontendPlugin_decompressed_Frontend_FETCH_FAULT_0 = FrontendPlugin_aligned_Frontend_FETCH_FAULT_0;
  assign FrontendPlugin_decompressed_Frontend_FETCH_FAULT_PAGE_0 = FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_0;
  assign FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_1 = FrontendPlugin_aligned_Frontend_INSTRUCTION_ALIGNED_1;
  assign FrontendPlugin_decompressed_Frontend_MASK_ALIGNED_1 = FrontendPlugin_aligned_Frontend_MASK_ALIGNED_1;
  assign FrontendPlugin_decompressed_PC_1 = FrontendPlugin_aligned_PC_1;
  assign FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_VALID_1 = FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1;
  assign FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_PC_NEXT_1 = FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_PC_NEXT_1;
  assign FrontendPlugin_decompressed_BRANCH_HISTORY_1 = FrontendPlugin_aligned_BRANCH_HISTORY_1;
  assign FrontendPlugin_decompressed_GSHARE_COUNTER_1_0 = FrontendPlugin_aligned_GSHARE_COUNTER_1_0;
  assign FrontendPlugin_decompressed_GSHARE_COUNTER_1_1 = FrontendPlugin_aligned_GSHARE_COUNTER_1_1;
  assign FrontendPlugin_decompressed_FETCH_ID_1 = FrontendPlugin_aligned_FETCH_ID_1;
  assign FrontendPlugin_decompressed_Frontend_FETCH_FAULT_1 = FrontendPlugin_aligned_Frontend_FETCH_FAULT_1;
  assign FrontendPlugin_decompressed_Frontend_FETCH_FAULT_PAGE_1 = FrontendPlugin_aligned_Frontend_FETCH_FAULT_PAGE_1;
  assign FrontendPlugin_decompressed_ready_output = FrontendPlugin_decoded_ready;
  assign FrontendPlugin_decoded_valid = FrontendPlugin_decompressed_valid;
  assign FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_0 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_DECOMPRESSED_0;
  assign FrontendPlugin_decoded_Frontend_INSTRUCTION_ALIGNED_0 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_0;
  assign FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_0 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_ILLEGAL_0;
  assign FrontendPlugin_decoded_Frontend_INSTRUCTION_DECOMPRESSED_1 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_DECOMPRESSED_1;
  assign FrontendPlugin_decoded_Frontend_INSTRUCTION_ALIGNED_1 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_ALIGNED_1;
  assign FrontendPlugin_decoded_Frontend_INSTRUCTION_ILLEGAL_1 = FrontendPlugin_decompressed_Frontend_INSTRUCTION_ILLEGAL_1;
  assign FrontendPlugin_decoded_Prediction_CONDITIONAL_TAKE_IT_0 = FrontendPlugin_decompressed_Prediction_CONDITIONAL_TAKE_IT_0;
  assign FrontendPlugin_decoded_GSHARE_COUNTER_0_0 = FrontendPlugin_decompressed_GSHARE_COUNTER_0_0;
  assign FrontendPlugin_decoded_GSHARE_COUNTER_0_1 = FrontendPlugin_decompressed_GSHARE_COUNTER_0_1;
  assign FrontendPlugin_decoded_Prediction_CONDITIONAL_TAKE_IT_1 = FrontendPlugin_decompressed_Prediction_CONDITIONAL_TAKE_IT_1;
  assign FrontendPlugin_decoded_GSHARE_COUNTER_1_0 = FrontendPlugin_decompressed_GSHARE_COUNTER_1_0;
  assign FrontendPlugin_decoded_GSHARE_COUNTER_1_1 = FrontendPlugin_decompressed_GSHARE_COUNTER_1_1;
  assign FrontendPlugin_decoded_FETCH_ID_0 = FrontendPlugin_decompressed_FETCH_ID_0;
  assign FrontendPlugin_decoded_FETCH_ID_1 = FrontendPlugin_decompressed_FETCH_ID_1;
  assign FrontendPlugin_decoded_Frontend_MASK_ALIGNED_0 = FrontendPlugin_decompressed_Frontend_MASK_ALIGNED_0;
  assign FrontendPlugin_decoded_Frontend_FETCH_FAULT_0 = FrontendPlugin_decompressed_Frontend_FETCH_FAULT_0;
  assign FrontendPlugin_decoded_Frontend_MASK_ALIGNED_1 = FrontendPlugin_decompressed_Frontend_MASK_ALIGNED_1;
  assign FrontendPlugin_decoded_Frontend_FETCH_FAULT_1 = FrontendPlugin_decompressed_Frontend_FETCH_FAULT_1;
  assign FrontendPlugin_decoded_Frontend_FETCH_FAULT_PAGE_0 = FrontendPlugin_decompressed_Frontend_FETCH_FAULT_PAGE_0;
  assign FrontendPlugin_decoded_Frontend_FETCH_FAULT_PAGE_1 = FrontendPlugin_decompressed_Frontend_FETCH_FAULT_PAGE_1;
  assign FrontendPlugin_decoded_PC_0 = FrontendPlugin_decompressed_PC_0;
  assign FrontendPlugin_decoded_PC_1 = FrontendPlugin_decompressed_PC_1;
  assign FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_0 = FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
  assign FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_1 = FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_PC_NEXT_1;
  assign FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_VALID_0 = FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_VALID_0;
  assign FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_VALID_1 = FrontendPlugin_decompressed_Prediction_ALIGNED_BRANCH_VALID_1;
  assign FrontendPlugin_decoded_BRANCH_HISTORY_0 = FrontendPlugin_decompressed_BRANCH_HISTORY_0;
  assign FrontendPlugin_decoded_BRANCH_HISTORY_1 = FrontendPlugin_decompressed_BRANCH_HISTORY_1;
  always @(*) begin
    FrontendPlugin_decoded_ready_output = FrontendPlugin_serialized_ready;
    if(when_Connection_l74_6) begin
      FrontendPlugin_decoded_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_6 = (! FrontendPlugin_serialized_valid);
  assign PcPlugin_logic_init_booted = PcPlugin_logic_init_counter[6];
  always @(*) begin
    PcPlugin_logic_fetchPc_correction = 1'b0;
    if(PcPlugin_logic_jump_pcLoad_valid) begin
      PcPlugin_logic_fetchPc_correction = 1'b1;
    end
  end

  assign PcPlugin_logic_fetchPc_output_fire = (PcPlugin_logic_fetchPc_output_valid && PcPlugin_logic_fetchPc_output_ready);
  assign PcPlugin_logic_fetchPc_corrected = (PcPlugin_logic_fetchPc_correction || PcPlugin_logic_fetchPc_correctionReg);
  assign PcPlugin_logic_fetchPc_pcRegPropagate = 1'b0;
  assign when_PcPlugin_l82 = (PcPlugin_logic_fetchPc_correction || PcPlugin_logic_fetchPc_pcRegPropagate);
  assign when_PcPlugin_l82_1 = ((! PcPlugin_logic_fetchPc_output_valid) && PcPlugin_logic_fetchPc_output_ready);
  always @(*) begin
    PcPlugin_logic_fetchPc_pc = (PcPlugin_logic_fetchPc_pcReg + _zz_PcPlugin_logic_fetchPc_pc);
    if(PcPlugin_logic_fetchPc_inc) begin
      PcPlugin_logic_fetchPc_pc[2 : 2] = 1'b0;
    end
    if(PcPlugin_logic_jump_pcLoad_valid) begin
      PcPlugin_logic_fetchPc_pc = PcPlugin_logic_jump_pcLoad_payload_pc;
    end
    PcPlugin_logic_fetchPc_pc[0] = 1'b0;
    PcPlugin_logic_fetchPc_pc[1] = 1'b0;
  end

  always @(*) begin
    PcPlugin_logic_fetchPc_flushed = 1'b0;
    if(PcPlugin_logic_jump_pcLoad_valid) begin
      PcPlugin_logic_fetchPc_flushed = 1'b1;
    end
  end

  assign when_PcPlugin_l98 = (PcPlugin_logic_init_booted && ((PcPlugin_logic_fetchPc_output_ready || PcPlugin_logic_fetchPc_correction) || PcPlugin_logic_fetchPc_pcRegPropagate));
  assign PcPlugin_logic_fetchPc_fetcherHalt = 1'b0;
  assign PcPlugin_logic_fetchPc_output_valid = ((! PcPlugin_logic_fetchPc_fetcherHalt) && PcPlugin_logic_init_booted);
  assign PcPlugin_logic_fetchPc_output_payload = PcPlugin_logic_fetchPc_pc;
  assign PcPlugin_logic_fetchPc_output_ready = FetchPlugin_stages_0_ready;
  assign FetchPlugin_stages_0_valid = PcPlugin_logic_fetchPc_output_valid;
  assign FetchPlugin_stages_0_Fetch_FETCH_PC = PcPlugin_logic_fetchPc_output_payload;
  always @(*) begin
    FetchPlugin_stages_1_Fetch_FETCH_PC_INC = (FetchPlugin_stages_1_Fetch_FETCH_PC + 32'h00000008);
    FetchPlugin_stages_1_Fetch_FETCH_PC_INC[2 : 0] = 3'b000;
  end

  assign fetchLastFire = FetchPlugin_stages_2_isFireing;
  assign fetchLastId = FetchPlugin_stages_2_FETCH_ID;
  assign AlignerPlugin_setup_s2m_isFlushed = FrontendPlugin_aligned_isFlushed;
  assign when_Connection_l66_1 = ({FrontendPlugin_aligned_isFlushed,_zz_FetchPlugin_stages_2_isFlushingRoot} != 2'b00);
  assign FetchPlugin_stages_2_isFlushed = when_Connection_l66_1;
  assign FetchPlugin_stages_1_isRemoved = (FetchPlugin_stages_1_isFlushed || FetchPlugin_stages_1_isThrown);
  assign when_Connection_l54 = ({when_Connection_l66_1,_zz_FetchPlugin_stages_1_isFlushingRoot} != 2'b00);
  assign FetchPlugin_stages_1_isFlushed = when_Connection_l54;
  assign FetchPlugin_stages_1_isFlushingNext = BtbPlugin_logic_applyIt_doIt;
  assign FetchPlugin_stages_1_isThrown = 1'b0;
  assign FetchPlugin_stages_0_isFlushed = (when_Connection_l54 || (BtbPlugin_logic_applyIt_doIt && 1'b1));
  assign FetchPlugin_stages_1_isFlushingRoot = (_zz_FetchPlugin_stages_1_isFlushingRoot != 1'b0);
  assign FetchPlugin_stages_2_isFlushingRoot = (_zz_FetchPlugin_stages_2_isFlushingRoot != 1'b0);
  assign AlignerPlugin_setup_s2m_isFlushingRoot = 1'b0;
  always @(*) begin
    _zz_FetchPlugin_stages_1_valid = FetchPlugin_stages_0_valid;
    if(when_Pipeline_l278_9) begin
      _zz_FetchPlugin_stages_1_valid = 1'b0;
    end
  end

  always @(*) begin
    FetchPlugin_stages_0_ready = FetchPlugin_stages_0_ready_output;
    if(when_Pipeline_l278_9) begin
      FetchPlugin_stages_0_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_9 = ({FetchPlugin_stages_0_haltRequest_MmuPlugin_l503,{FetchPlugin_stages_0_haltRequest_PrivilegedPlugin_l968,{FetchPlugin_stages_0_haltRequest_Lsu2Plugin_l1548,{FetchPlugin_stages_0_haltRequest_EnvCallPlugin_l125,{FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l583,{FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l552,{FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l476,FetchPlugin_stages_0_haltRequest_FetchCachePlugin_l389}}}}}}} != 8'h00);
  always @(*) begin
    _zz_FetchPlugin_stages_2_valid = FetchPlugin_stages_1_valid;
    if(FetchPlugin_stages_1_isFlushingRoot) begin
      _zz_FetchPlugin_stages_2_valid = 1'b0;
    end
  end

  assign FetchPlugin_stages_1_ready = FetchPlugin_stages_1_ready_output;
  always @(*) begin
    _zz_AlignerPlugin_setup_s2m_valid = FetchPlugin_stages_2_valid;
    if(FetchPlugin_stages_2_isFlushingRoot) begin
      _zz_AlignerPlugin_setup_s2m_valid = 1'b0;
    end
  end

  assign FetchPlugin_stages_2_ready = FetchPlugin_stages_2_ready_output;
  always @(*) begin
    AlignerPlugin_setup_s2m_ready = 1'b1;
    if(when_Pipeline_l278_10) begin
      AlignerPlugin_setup_s2m_ready = 1'b0;
    end
  end

  assign when_Pipeline_l278_10 = (AlignerPlugin_setup_s2m_haltRequest_AlignerPlugin_l270 != 1'b0);
  always @(*) begin
    FetchPlugin_stages_0_ready_output = FetchPlugin_stages_1_ready;
    if(when_Connection_l74_7) begin
      FetchPlugin_stages_0_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_7 = (! FetchPlugin_stages_1_valid);
  always @(*) begin
    FetchPlugin_stages_1_ready_output = FetchPlugin_stages_2_ready;
    if(when_Connection_l74_8) begin
      FetchPlugin_stages_1_ready_output = 1'b1;
    end
  end

  assign when_Connection_l74_8 = (! FetchPlugin_stages_2_valid);
  assign FetchPlugin_stages_2_ready_output = (! FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid);
  assign AlignerPlugin_setup_s2m_valid = (_zz_AlignerPlugin_setup_s2m_valid || FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid);
  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_WORD = FetchPlugin_stages_2_Fetch_WORD_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_WORD = FetchPlugin_stages_2_Fetch_WORD;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_FETCH_PC = FetchPlugin_stages_2_Fetch_FETCH_PC_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_FETCH_PC = FetchPlugin_stages_2_Fetch_FETCH_PC;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_WORD_FAULT = FetchPlugin_stages_2_Fetch_WORD_FAULT_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_WORD_FAULT = FetchPlugin_stages_2_Fetch_WORD_FAULT;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE = FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE = FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_BRANCH_HISTORY = FetchPlugin_stages_2_BRANCH_HISTORY_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_BRANCH_HISTORY = FetchPlugin_stages_2_BRANCH_HISTORY;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_FETCH_ID = FetchPlugin_stages_2_FETCH_ID_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_FETCH_ID = FetchPlugin_stages_2_FETCH_ID;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_SLICE = FetchPlugin_stages_2_Prediction_WORD_BRANCH_SLICE_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_SLICE = FetchPlugin_stages_2_Prediction_WORD_BRANCH_SLICE;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID = FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID = FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_MASK_FRONT = FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_MASK_FRONT = FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT = FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT = FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_SLICE = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_SLICE_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_SLICE = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_SLICE;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE = FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_GSHARE_COUNTER_0 = FetchPlugin_stages_2_GSHARE_COUNTER_s2mBuffer_0;
    end else begin
      AlignerPlugin_setup_s2m_GSHARE_COUNTER_0 = FetchPlugin_stages_2_GSHARE_COUNTER_0;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_GSHARE_COUNTER_1 = FetchPlugin_stages_2_GSHARE_COUNTER_s2mBuffer_1;
    end else begin
      AlignerPlugin_setup_s2m_GSHARE_COUNTER_1 = FetchPlugin_stages_2_GSHARE_COUNTER_1;
    end
  end

  always @(*) begin
    if(FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid) begin
      AlignerPlugin_setup_s2m_Fetch_FETCH_PC_INC = FetchPlugin_stages_2_Fetch_FETCH_PC_INC_s2mBuffer;
    end else begin
      AlignerPlugin_setup_s2m_Fetch_FETCH_PC_INC = FetchPlugin_stages_2_Fetch_FETCH_PC_INC;
    end
  end

  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_stateReg;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
        if(PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW;
        end else begin
          if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
            PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW;
          end else begin
            if(PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid) begin
              PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE;
            end
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
        if(PerformanceCounterPlugin_setup_readPort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH;
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
        if(PerformanceCounterPlugin_logic_fsm_cmd_flusher) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW;
        end else begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_IDLE;
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
        if(PerformanceCounterPlugin_setup_writePort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH;
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
        if(PerformanceCounterPlugin_setup_readPort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_CALC;
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
        if(PerformanceCounterPlugin_setup_writePort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_IDLE;
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
        if(PerformanceCounterPlugin_setup_writePort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION;
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
        PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_IDLE;
      end
      default : begin
      end
    endcase
    if(PerformanceCounterPlugin_logic_fsm_wantStart) begin
      PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_IDLE;
    end
    if(PerformanceCounterPlugin_logic_fsm_wantKill) begin
      PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_enumDef_BOOT;
    end
  end

  assign when_PerformanceCounterPlugin_l201 = PerformanceCounterPlugin_logic_fsm_counterReaded[5];
  assign when_PerformanceCounterPlugin_l161 = (! PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_high);
  assign when_PerformanceCounterPlugin_l169 = (PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address == 3'b010);
  always @(*) begin
    PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_stateReg;
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
        if(PrivilegedPlugin_logic_rescheduleUnbuffered_valid) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_SETUP;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
        if(when_PrivilegedPlugin_l766) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ;
        end else begin
          case(PrivilegedPlugin_logic_reschedule_payload_cause)
            4'b1001 : begin
              PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC;
            end
            4'b1010 : begin
              PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC;
            end
            4'b1000 : begin
              PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_EPC_READ;
            end
            default : begin
              PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ;
            end
          endcase
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        if(PrivilegedPlugin_setup_ramWrite_ready) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_TRAP;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        if(PrivilegedPlugin_setup_ramWrite_ready) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        if(PrivilegedPlugin_setup_ramRead_ready) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_XRET;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        if(PrivilegedPlugin_setup_ramRead_ready) begin
          PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE;
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
        PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_IDLE;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
        PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
        PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_IDLE;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
        PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_IDLE;
      end
      default : begin
      end
    endcase
    if(PrivilegedPlugin_logic_fsm_wantStart) begin
      PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_IDLE;
    end
    if(PrivilegedPlugin_logic_fsm_wantKill) begin
      PrivilegedPlugin_logic_fsm_stateNext = PrivilegedPlugin_logic_fsm_enumDef_BOOT;
    end
  end

  assign when_PrivilegedPlugin_l766 = ((! PrivilegedPlugin_logic_reschedule_payload_fromCommit) && PrivilegedPlugin_logic_decoderInterrupt_raised);
  always @(*) begin
    _zz_PrivilegedPlugin_setup_ramWrite_address = 5'h15;
    case(PrivilegedPlugin_logic_fsm_trap_targetPrivilege)
      2'b01 : begin
        _zz_PrivilegedPlugin_setup_ramWrite_address = 5'h11;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_PrivilegedPlugin_setup_ramWrite_address_1 = 5'h16;
    case(PrivilegedPlugin_logic_fsm_trap_targetPrivilege)
      2'b01 : begin
        _zz_PrivilegedPlugin_setup_ramWrite_address_1 = 5'h12;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_PrivilegedPlugin_setup_ramRead_address = 5'h15;
    case(PrivilegedPlugin_logic_fsm_xret_sourcePrivilege)
      2'b01 : begin
        _zz_PrivilegedPlugin_setup_ramRead_address = 5'h11;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_PrivilegedPlugin_setup_ramRead_address_1 = 5'h17;
    case(PrivilegedPlugin_logic_fsm_trap_targetPrivilege)
      2'b01 : begin
        _zz_PrivilegedPlugin_setup_ramRead_address_1 = 5'h13;
      end
      default : begin
      end
    endcase
  end

  assign when_PrivilegedPlugin_l952 = (PrivilegedPlugin_logic_fsm_xret_targetPrivilege < 2'b11);
  assign switch_PrivilegedPlugin_l953 = PrivilegedPlugin_logic_reschedule_payload_tval[1 : 0];
  assign when_StateMachine_l253_2 = ((! (PrivilegedPlugin_logic_fsm_stateReg == PrivilegedPlugin_logic_fsm_enumDef_IDLE)) && (PrivilegedPlugin_logic_fsm_stateNext == PrivilegedPlugin_logic_fsm_enumDef_IDLE));
  always @(*) begin
    _zz_FetchCachePlugin_logic_banks_0_read_rsp = _zz_FetchCachePlugin_logic_banks_0_mem_port1;
    if(when_MultiportRam_l328) begin
      _zz_FetchCachePlugin_logic_banks_0_read_rsp = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    _zz_FetchCachePlugin_logic_banks_1_read_rsp = _zz_FetchCachePlugin_logic_banks_1_mem_port1;
    if(when_MultiportRam_l328_1) begin
      _zz_FetchCachePlugin_logic_banks_1_read_rsp = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    _zz_FetchCachePlugin_logic_banks_2_read_rsp = _zz_FetchCachePlugin_logic_banks_2_mem_port1;
    if(when_MultiportRam_l328_2) begin
      _zz_FetchCachePlugin_logic_banks_2_read_rsp = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    _zz_FetchCachePlugin_logic_banks_3_read_rsp = _zz_FetchCachePlugin_logic_banks_3_mem_port1;
    if(when_MultiportRam_l328_3) begin
      _zz_FetchCachePlugin_logic_banks_3_read_rsp = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(*) begin
    _zz_FetchPlugin_stages_1_GSHARE_COUNTER_0_1 = _zz_GSharePlugin_logic_mem_counter_port1;
    if(when_MultiportRam_l328_4) begin
      _zz_FetchPlugin_stages_1_GSHARE_COUNTER_0_1 = 4'bxxxx;
    end
  end

  always @(*) begin
    _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_2 = _zz_Lsu2Plugin_logic_lq_hazardPrediction_mem_port1;
    if(when_MultiportRam_l362) begin
      _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_2 = _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_3;
    end
  end

  always @(*) begin
    _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter_1 = _zz_Lsu2Plugin_logic_lq_hitPrediction_mem_port1;
    if(when_MultiportRam_l362_1) begin
      _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter_1 = _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter_2;
    end
  end

  assign BranchContextPlugin_logic_mem_earlyBranch_io_writes_0_payload_data = {FrontendPlugin_allocated_BRANCH_EARLY_0_pc,FrontendPlugin_allocated_BRANCH_EARLY_0_taken};
  assign BranchContextPlugin_logic_mem_earlyBranch_io_writes_1_payload_data = {FrontendPlugin_allocated_BRANCH_EARLY_1_pc,FrontendPlugin_allocated_BRANCH_EARLY_1_taken};
  assign BranchContextPlugin_logic_mem_earlyBranch_io_read_0_cmd_valid = 1'b1;
  assign BranchContextPlugin_logic_mem_earlyBranch_io_read_1_cmd_valid = 1'b1;
  assign BranchContextPlugin_logic_mem_finalBranch_io_writes_0_payload_data = {ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_taken,{ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcTarget,ALU0_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice}};
  assign BranchContextPlugin_logic_mem_finalBranch_io_writes_1_payload_data = {ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_taken,{ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcTarget,ALU1_BranchPlugin_logic_branch_finalBranch_payload_data_pcOnLastSlice}};
  assign BranchContextPlugin_logic_mem_finalBranch_io_read_0_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_io_writes_0_payload_data = Lsu2Plugin_logic_allocation_stores_alloc;
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_io_writes_1_payload_data = Lsu2Plugin_logic_allocation_stores_alloc_1;
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_0_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_1_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_1_cmd_payload = AguPlugin_setup_port_payload_aguId[3:0];
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_2_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_lq_mem_sqAlloc_io_read_3_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_lq_mem_doSpecial_io_writes_0_payload_data = 1'b0;
  assign Lsu2Plugin_logic_lq_mem_doSpecial_io_writes_1_payload_data = 1'b0;
  assign Lsu2Plugin_logic_lq_mem_doSpecial_io_writes_2_payload_data = 1'b1;
  assign Lsu2Plugin_logic_lq_mem_doSpecial_io_read_0_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_lq_mem_needTranslation_io_writes_0_payload_address = AguPlugin_setup_port_payload_aguId[3:0];
  assign Lsu2Plugin_logic_lq_mem_needTranslation_io_writes_0_payload_data = 1'b1;
  assign Lsu2Plugin_logic_lq_mem_needTranslation_io_writes_1_payload_data = Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO;
  assign Lsu2Plugin_logic_lq_mem_needTranslation_io_read_0_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_sq_mem_needTranslation_io_writes_0_payload_address = AguPlugin_setup_port_payload_aguId[3:0];
  assign Lsu2Plugin_logic_sq_mem_needTranslation_io_writes_0_payload_data = 1'b1;
  assign Lsu2Plugin_logic_sq_mem_needTranslation_io_writes_1_payload_data = Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO;
  assign Lsu2Plugin_logic_sq_mem_needTranslation_io_read_0_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_sq_mem_needTranslation_io_read_1_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_sq_mem_feededOnce_io_writes_0_payload_data = 1'b0;
  assign Lsu2Plugin_logic_sq_mem_feededOnce_io_writes_1_payload_data = 1'b0;
  assign Lsu2Plugin_logic_sq_mem_feededOnce_io_writes_2_payload_data = 1'b1;
  assign Lsu2Plugin_logic_sq_mem_feededOnce_io_read_0_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_sq_mem_doSpecial_io_writes_0_payload_data = 1'b0;
  assign Lsu2Plugin_logic_sq_mem_doSpecial_io_writes_1_payload_data = 1'b0;
  assign Lsu2Plugin_logic_sq_mem_doSpecial_io_writes_2_payload_data = 1'b1;
  assign Lsu2Plugin_logic_sq_mem_doSpecial_io_read_0_cmd_valid = 1'b1;
  assign Lsu2Plugin_logic_sq_mem_lqAlloc_io_writes_0_payload_data = Lsu2Plugin_logic_allocation_loads_alloc_1;
  assign Lsu2Plugin_logic_sq_mem_lqAlloc_io_writes_1_payload_data = Lsu2Plugin_logic_allocation_loads_alloc_2;
  assign Lsu2Plugin_logic_sq_mem_lqAlloc_io_read_0_cmd_valid = 1'b1;
  assign BranchContextPlugin_free_dispatchMem_mem_io_read_0_cmd_valid = 1'b1;
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_0_valid = (ALU0_ExecutionUnitBase_pipeline_execute_1_isFireing && 1'b1);
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_0_payload_data = ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND;
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_1_valid = (ALU1_ExecutionUnitBase_pipeline_execute_1_isFireing && 1'b1);
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_writes_1_payload_data = ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND;
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_0_cmd_valid = 1'b1;
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_0_cmd_payload = {_zz_io_read_0_cmd_payload,1'b0};
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_1_cmd_valid = 1'b1;
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_1_cmd_payload = {_zz_io_read_0_cmd_payload,1'b1};
  assign RobPlugin_logic_storage_BRANCH_TAKEN_banks_0_io_read_2_cmd_valid = 1'b1;
  assign CommitPlugin_logic_free_lineEventStream_fifo_io_flush = 1'b0;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      HistoryPlugin_logic_update_pushes_2_state <= 24'h000000;
      HistoryPlugin_logic_update_pushes_0_state <= 24'h000000;
      PrivilegedPlugin_setup_privilege <= 2'b11;
      FetchPlugin_stages_1_FETCH_ID <= 12'h000;
      _zz_FetchPlugin_stages_1_isFirstCycle <= 1'b0;
      FetchCachePlugin_logic_invalidate_requested <= 1'b0;
      FetchCachePlugin_logic_invalidate_counter <= 7'h00;
      FetchCachePlugin_logic_invalidate_firstEver <= 1'b1;
      FetchCachePlugin_logic_invalidate_done_regNext <= 1'b0;
      FetchCachePlugin_logic_refill_valid <= 1'b0;
      FetchCachePlugin_logic_refill_hadError <= 1'b0;
      FetchCachePlugin_logic_refill_pushCounter <= 32'h00000000;
      FetchCachePlugin_logic_refill_cmdSent <= 1'b0;
      FetchCachePlugin_logic_refill_randomWay_value <= 2'b00;
      FetchCachePlugin_logic_refill_wordIndex <= 3'b000;
      FetchCachePlugin_logic_refill_fire_regNext <= 1'b0;
      AlignerPlugin_logic_buffer_mask <= 2'b00;
      AlignerPlugin_logic_correctionSent <= 1'b0;
      DispatchPlugin_logic_sparseRob_todo <= 2'b11;
      BranchContextPlugin_logic_ptr_alloc <= 5'h00;
      BranchContextPlugin_logic_ptr_commited <= 5'h00;
      BranchContextPlugin_logic_ptr_free <= 5'h00;
      HistoryPlugin_logic_onCommit_value <= 24'h000000;
      DecoderPredictionPlugin_logic_ras_ptr_push <= 4'b0000;
      DecoderPredictionPlugin_logic_ras_ptr_pop <= 4'b1111;
      BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      toplevel_DataCachePlugin_logic_cache_io_refillEvent_regNext <= 1'b0;
      toplevel_DataCachePlugin_logic_cache_io_writebackEvent_regNext <= 1'b0;
      _zz_DataCachePlugin_logic_load_ohHistory_1 <= 2'b00;
      _zz_DataCachePlugin_logic_load_ohHistory_2 <= 2'b00;
      CommitPlugin_logic_ptr_alloc <= 7'h00;
      CommitPlugin_logic_ptr_commit <= 7'h00;
      CommitPlugin_logic_ptr_free <= 7'h00;
      CommitPlugin_logic_ptr_empty <= 1'b1;
      CommitPlugin_logic_reschedule_fresh <= 1'b0;
      CommitPlugin_logic_reschedule_valid <= 1'b0;
      CommitPlugin_logic_commit_mask <= 2'b11;
      CommitDebugFilterPlugin_logic_filters_0_value <= 32'h00000000;
      CommitDebugFilterPlugin_logic_filters_1_value <= 32'h00000000;
      CommitDebugFilterPlugin_logic_filters_2_value <= 32'h00000000;
      PrivilegedPlugin_logic_machine_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_machine_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_machine_mstatus_mie <= 1'b0;
      PrivilegedPlugin_logic_machine_mstatus_mpie <= 1'b0;
      PrivilegedPlugin_logic_machine_mstatus_mpp <= 2'b00;
      PrivilegedPlugin_logic_machine_mstatus_fs <= 2'b00;
      PrivilegedPlugin_logic_machine_mip_meip <= 1'b0;
      PrivilegedPlugin_logic_machine_mip_mtip <= 1'b0;
      PrivilegedPlugin_logic_machine_mip_msip <= 1'b0;
      PrivilegedPlugin_logic_machine_mie_meie <= 1'b0;
      PrivilegedPlugin_logic_machine_mie_mtie <= 1'b0;
      PrivilegedPlugin_logic_machine_mie_msie <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_iam <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_bp <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_eu <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_es <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_ipf <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_lpf <= 1'b0;
      PrivilegedPlugin_logic_machine_medeleg_spf <= 1'b0;
      PrivilegedPlugin_logic_machine_mideleg_st <= 1'b0;
      PrivilegedPlugin_logic_machine_mideleg_se <= 1'b0;
      PrivilegedPlugin_logic_machine_mideleg_ss <= 1'b0;
      PrivilegedPlugin_logic_supervisor_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_supervisor_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_supervisor_sstatus_sie <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sstatus_spie <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sstatus_spp <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sip_seipSoft <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sip_stip <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sip_ssip <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sie_seie <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sie_stie <= 1'b0;
      PrivilegedPlugin_logic_supervisor_sie_ssie <= 1'b0;
      PrivilegedPlugin_logic_rescheduleUnbuffered_rValid <= 1'b0;
      _zz_PerformanceCounterPlugin_logic_branchMissEvent <= 1'b0;
      PerformanceCounterPlugin_logic_ignoreNextCommit <= 1'b0;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded <= 6'h00;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2 <= 6'h00;
      PerformanceCounterPlugin_logic_commitCount_regNext <= 2'b00;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3 <= 6'h00;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4 <= 6'h00;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5 <= 6'h00;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6 <= 6'h00;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_7 <= 3'b000;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_8 <= 3'b000;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_9 <= 3'b000;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_10 <= 3'b000;
      EU0_DivPlugin_logic_feed_cmdSent <= 1'b0;
      AguPlugin_logic_fired <= 1'b0;
      EnvCallPlugin_logic_flushes_stateReg <= EnvCallPlugin_logic_flushes_enumDef_BOOT;
      integer_RfTranslationPlugin_logic_init_counter <= 6'h00;
      integer_RfAllocationPlugin_logic_init_counter <= 7'h01;
      HistoryPlugin_logic_onFetch_value <= 24'h000000;
      Lsu2Plugin_logic_lq_regs_0_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_8_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_8_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_8_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_9_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_9_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_9_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_10_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_10_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_10_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_11_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_11_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_11_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_12_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_12_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_12_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_13_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_13_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_13_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_14_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_14_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_14_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_regs_15_valid <= 1'b0;
      Lsu2Plugin_logic_lq_regs_15_redo <= 1'b0;
      Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefill <= 2'b00;
      Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_lq_regs_15_waitOn_sqWriteback <= 1'b0;
      Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeed <= 1'b0;
      Lsu2Plugin_logic_lq_ptr_priority <= 15'h0000;
      Lsu2Plugin_logic_lq_ptr_alloc <= 5'h00;
      Lsu2Plugin_logic_lq_ptr_free <= 5'h00;
      Lsu2Plugin_logic_lq_tracker_free <= 5'h10;
      Lsu2Plugin_logic_lq_reservation_valid <= 1'b0;
      Lsu2Plugin_logic_lq_reservation_counter <= 7'h00;
      Lsu2Plugin_logic_sq_regs_0_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_0_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_0_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_1_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_1_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_1_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_2_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_2_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_2_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_3_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_3_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_3_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_4_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_4_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_4_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_5_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_5_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_5_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_6_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_6_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_6_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_7_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_7_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_7_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_8_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_8_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_8_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_9_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_9_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_9_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_10_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_10_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_10_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_11_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_11_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_11_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_12_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_12_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_12_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_13_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_13_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_13_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_14_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_14_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_14_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_regs_15_valid <= 1'b0;
      Lsu2Plugin_logic_sq_regs_15_redo <= 1'b0;
      Lsu2Plugin_logic_sq_regs_15_commited <= 1'b0;
      Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAny <= 1'b0;
      Lsu2Plugin_logic_sq_ptr_priority <= 15'h0000;
      Lsu2Plugin_logic_sq_ptr_alloc <= 5'h00;
      Lsu2Plugin_logic_sq_ptr_commit <= 5'h00;
      Lsu2Plugin_logic_sq_ptr_writeBack <= 5'h00;
      Lsu2Plugin_logic_sq_ptr_free <= 5'h00;
      Lsu2Plugin_logic_sq_ptr_onFreeLast_valid <= 1'b0;
      Lsu2Plugin_logic_sq_tracker_free <= 5'h10;
      Lsu2Plugin_logic_sharedPip_speculativeHitPredictionGotReschedule <= 1'b0;
      Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled <= 1'b1;
      Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask <= 1'b1;
      Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask <= 1'b1;
      Lsu2Plugin_logic_writeback_generation <= 1'b0;
      Lsu2Plugin_logic_writeback_waitOn_refillSlot <= 2'b00;
      Lsu2Plugin_logic_writeback_waitOn_refillSlotAny <= 1'b0;
      toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rValid <= 1'b0;
      Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_valid <= 1'b0;
      Lsu2Plugin_logic_flush_busy <= 1'b0;
      Lsu2Plugin_logic_flush_doit <= 1'b0;
      LsuPlugin_peripheralBus_rsp_valid_regNext <= 1'b0;
      Lsu2Plugin_logic_special_enabled <= 1'b0;
      Lsu2Plugin_logic_special_cmdSent <= 1'b0;
      Lsu2Plugin_logic_special_atomic_lockDelayCounter <= 2'b00;
      Lsu2Plugin_logic_special_atomic_comp_wakeRf <= 1'b0;
      Lsu2Plugin_logic_special_atomic_comp_rfWrite <= 1'b0;
      MmuPlugin_logic_satp_mode <= 1'b0;
      MmuPlugin_logic_satp_ppn <= 20'h00000;
      MmuPlugin_logic_status_mxr <= 1'b0;
      MmuPlugin_logic_status_sum <= 1'b0;
      MmuPlugin_logic_status_mprv <= 1'b0;
      FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value <= 2'b00;
      FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value <= 1'b0;
      Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value <= 2'b00;
      Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value <= 1'b0;
      Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg <= 1'b1;
      Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg <= 1'b1;
      PrivilegedPlugin_logic_decoderInterrupt_raised <= 1'b0;
      PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt <= 1'b0;
      PrivilegedPlugin_logic_decoderInterrupt_counter <= 3'b000;
      PerformanceCounterPlugin_logic_fsm_done <= 1'b0;
      PerformanceCounterPlugin_logic_csrRead_fired <= 1'b0;
      PerformanceCounterPlugin_logic_csrWrite_fired <= 1'b0;
      FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg <= 1'b1;
      MmuPlugin_logic_refill_cacheRefill <= 2'b00;
      MmuPlugin_logic_refill_cacheRefillAny <= 1'b0;
      MmuPlugin_logic_refill_load_rsp_valid <= 1'b0;
      MmuPlugin_logic_invalidate_requested <= 1'b1;
      MmuPlugin_logic_invalidate_counter <= 6'h00;
      MmuPlugin_logic_invalidate_done_regNext <= 1'b0;
      Lsu2Plugin_logic_sharedPip_stages_1_valid <= 1'b0;
      Lsu2Plugin_logic_sharedPip_stages_2_valid <= 1'b0;
      Lsu2Plugin_logic_sharedPip_stages_3_valid <= 1'b0;
      Lsu2Plugin_logic_lqSqArbitration_s1_valid <= 1'b0;
      Lsu2Plugin_logic_special_atomic_stateReg <= Lsu2Plugin_logic_special_atomic_enumDef_BOOT;
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_enumDef_BOOT;
      CsrRamPlugin_logic_flush_counter <= 6'h00;
      EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired <= 1'b0;
      EU0_CsrAccessPlugin_logic_fsm_stateReg <= EU0_CsrAccessPlugin_logic_fsm_enumDef_BOOT;
      DecoderPlugin_logic_exception_trigged <= 1'b0;
      DecoderPlugin_logic_exception_doItAgain <= 1'b0;
      FrontendPlugin_decoded_OP_ID <= 12'h000;
      DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle <= 1'b1;
      ALU0_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      ALU0_ExecutionUnitBase_pipeline_execute_1_valid <= 1'b0;
      ALU1_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      ALU1_ExecutionUnitBase_pipeline_execute_1_valid <= 1'b0;
      EU0_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      EU0_ExecutionUnitBase_pipeline_execute_1_valid <= 1'b0;
      EU0_ExecutionUnitBase_pipeline_execute_2_valid <= 1'b0;
      DispatchPlugin_logic_ptr_next <= 6'h22;
      DispatchPlugin_logic_ptr_current <= 6'h20;
      DispatchPlugin_logic_push_fenceYoungerLast <= 1'b0;
      DispatchPlugin_logic_pop_0_stagesList_1_valid <= 1'b0;
      DispatchPlugin_logic_pop_1_stagesList_1_valid <= 1'b0;
      DispatchPlugin_logic_pop_2_stagesList_1_valid <= 1'b0;
      RfDependencyPlugin_logic_forRf_integer_init_counter <= 7'h00;
      FrontendPlugin_dispatch_valid <= 1'b0;
      FrontendPlugin_serialized_valid <= 1'b0;
      PcPlugin_logic_init_counter <= 7'h00;
      PcPlugin_logic_fetchPc_pcReg <= 32'h80000000;
      PcPlugin_logic_fetchPc_correctionReg <= 1'b0;
      PcPlugin_logic_fetchPc_inc <= 1'b0;
      FetchPlugin_stages_1_valid <= 1'b0;
      FetchPlugin_stages_2_valid <= 1'b0;
      FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid <= 1'b0;
      PerformanceCounterPlugin_logic_fsm_stateReg <= PerformanceCounterPlugin_logic_fsm_enumDef_BOOT;
      PrivilegedPlugin_logic_fsm_stateReg <= PrivilegedPlugin_logic_fsm_enumDef_BOOT;
      when_MultiportRam_l328 <= 1'b0;
      when_MultiportRam_l328_1 <= 1'b0;
      when_MultiportRam_l328_2 <= 1'b0;
      when_MultiportRam_l328_3 <= 1'b0;
      when_MultiportRam_l328_4 <= 1'b0;
      when_MultiportRam_l362 <= 1'b0;
      when_MultiportRam_l362_1 <= 1'b0;
    end else begin
      FetchPlugin_stages_1_FETCH_ID <= (FetchPlugin_stages_1_FETCH_ID + _zz_FetchPlugin_stages_1_FETCH_ID);
      if(FetchPlugin_stages_1_valid) begin
        _zz_FetchPlugin_stages_1_isFirstCycle <= 1'b1;
      end
      if(when_Stage_l170) begin
        _zz_FetchPlugin_stages_1_isFirstCycle <= 1'b0;
      end
      if(FetchCachePlugin_setup_invalidatePort_cmd_valid) begin
        FetchCachePlugin_logic_invalidate_requested <= 1'b1;
      end
      if(FetchCachePlugin_logic_invalidate_done) begin
        FetchCachePlugin_logic_invalidate_firstEver <= 1'b0;
      end
      if(when_FetchCachePlugin_l379) begin
        FetchCachePlugin_logic_invalidate_counter <= (FetchCachePlugin_logic_invalidate_counter + 7'h01);
      end
      if(when_FetchCachePlugin_l391) begin
        FetchCachePlugin_logic_invalidate_counter <= 7'h00;
        FetchCachePlugin_logic_invalidate_requested <= 1'b0;
      end
      FetchCachePlugin_logic_invalidate_done_regNext <= FetchCachePlugin_logic_invalidate_done;
      if(FetchCachePlugin_logic_refill_fire) begin
        FetchCachePlugin_logic_refill_valid <= 1'b0;
      end
      if(when_FetchCachePlugin_l422) begin
        if(FetchCachePlugin_logic_refill_start_valid) begin
          FetchCachePlugin_logic_refill_valid <= 1'b1;
          FetchCachePlugin_logic_refill_pushCounter <= (FetchCachePlugin_logic_refill_pushCounter + 32'h00000001);
        end
      end
      if(FetchCachePlugin_mem_cmd_fire) begin
        FetchCachePlugin_logic_refill_cmdSent <= 1'b1;
      end
      if(FetchCachePlugin_logic_refill_fire) begin
        FetchCachePlugin_logic_refill_cmdSent <= 1'b0;
      end
      FetchCachePlugin_logic_refill_randomWay_value <= FetchCachePlugin_logic_refill_randomWay_valueNext;
      if(FetchCachePlugin_mem_rsp_valid) begin
        FetchCachePlugin_logic_refill_wordIndex <= (FetchCachePlugin_logic_refill_wordIndex + 3'b001);
        if(FetchCachePlugin_mem_rsp_payload_error) begin
          FetchCachePlugin_logic_refill_hadError <= 1'b1;
        end
      end
      if(FetchCachePlugin_logic_refill_fire) begin
        FetchCachePlugin_logic_refill_hadError <= 1'b0;
      end
      FetchCachePlugin_logic_refill_fire_regNext <= FetchCachePlugin_logic_refill_fire;
      if(AlignerPlugin_logic_fireOutput) begin
        AlignerPlugin_logic_buffer_mask <= AlignerPlugin_logic_slices_remains_2[1 : 0];
      end
      if(AlignerPlugin_logic_fireInput) begin
        AlignerPlugin_logic_buffer_mask <= ((AlignerPlugin_logic_fireOutput ? AlignerPlugin_logic_slices_remains_2[3 : 2] : AlignerPlugin_setup_s2m_MASK_FRONT) & AlignerPlugin_logic_postMask);
      end
      if(AlignerPlugin_setup_sequenceJump_valid) begin
        AlignerPlugin_logic_correctionSent <= 1'b1;
      end
      if(when_AlignerPlugin_l264) begin
        AlignerPlugin_logic_correctionSent <= 1'b0;
      end
      if(FrontendPlugin_aligned_isFlushed) begin
        AlignerPlugin_logic_buffer_mask <= 2'b00;
      end
      if(FrontendPlugin_serialized_isForked) begin
        DispatchPlugin_logic_sparseRob_todo <= (DispatchPlugin_logic_sparseRob_todo & (~ DispatchPlugin_logic_sparseRob_filter));
      end
      if(when_DispatchPlugin_l94) begin
        DispatchPlugin_logic_sparseRob_todo <= 2'b11;
      end
      if(FrontendPlugin_allocated_isFireing) begin
        BranchContextPlugin_logic_ptr_alloc <= BranchContextPlugin_logic_alloc_allocNext_2;
      end
      DecoderPredictionPlugin_logic_ras_ptr_push <= (_zz_DecoderPredictionPlugin_logic_ras_ptr_push - _zz_DecoderPredictionPlugin_logic_ras_ptr_push_3);
      DecoderPredictionPlugin_logic_ras_ptr_pop <= (_zz_DecoderPredictionPlugin_logic_ras_ptr_pop - _zz_DecoderPredictionPlugin_logic_ras_ptr_pop_3);
      if(FetchPlugin_stages_1_valid) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b1;
      end
      if(when_BtbPlugin_l109) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      end
      toplevel_DataCachePlugin_logic_cache_io_refillEvent_regNext <= DataCachePlugin_logic_cache_io_refillEvent;
      toplevel_DataCachePlugin_logic_cache_io_writebackEvent_regNext <= DataCachePlugin_logic_cache_io_writebackEvent;
      _zz_DataCachePlugin_logic_load_ohHistory_1 <= _zz_DataCachePlugin_logic_load_ohHistory_0;
      _zz_DataCachePlugin_logic_load_ohHistory_2 <= _zz_DataCachePlugin_logic_load_ohHistory_1;
      CommitPlugin_logic_ptr_commit <= CommitPlugin_logic_ptr_commitNext;
      CommitPlugin_logic_ptr_alloc <= CommitPlugin_logic_ptr_allocNext;
      CommitPlugin_logic_ptr_empty <= (CommitPlugin_logic_ptr_allocNext == CommitPlugin_logic_ptr_commitNext);
      CommitPlugin_logic_reschedule_fresh <= 1'b0;
      if(when_CommitPlugin_l131) begin
        CommitPlugin_logic_reschedule_fresh <= 1'b1;
        CommitPlugin_logic_reschedule_valid <= 1'b1;
      end
      CommitPlugin_logic_commit_mask <= CommitPlugin_logic_commit_maskComb;
      if(CommitPlugin_logic_commit_rescheduleHit) begin
        CommitPlugin_logic_reschedule_valid <= 1'b0;
      end
      if(when_CommitPlugin_l194) begin
        if(when_CommitPlugin_l217) begin
          CommitPlugin_logic_commit_mask <= 2'b11;
        end
      end
      if(CommitPlugin_logic_ptr_canFree) begin
        CommitPlugin_logic_ptr_free <= (CommitPlugin_logic_ptr_free + 7'h02);
      end
      CommitDebugFilterPlugin_logic_filters_0_value <= (CommitDebugFilterPlugin_logic_filters_0_value + _zz_CommitDebugFilterPlugin_logic_filters_0_value);
      CommitDebugFilterPlugin_logic_filters_1_value <= (CommitDebugFilterPlugin_logic_filters_1_value + _zz_CommitDebugFilterPlugin_logic_filters_1_value);
      CommitDebugFilterPlugin_logic_filters_2_value <= (CommitDebugFilterPlugin_logic_filters_2_value + _zz_CommitDebugFilterPlugin_logic_filters_2_value);
      PrivilegedPlugin_logic_machine_mip_meip <= PrivilegedPlugin_io_int_machine_external;
      PrivilegedPlugin_logic_machine_mip_mtip <= PrivilegedPlugin_io_int_machine_timer;
      PrivilegedPlugin_logic_machine_mip_msip <= PrivilegedPlugin_io_int_machine_software;
      if(PrivilegedPlugin_logic_rescheduleUnbuffered_ready) begin
        PrivilegedPlugin_logic_rescheduleUnbuffered_rValid <= PrivilegedPlugin_logic_rescheduleUnbuffered_valid;
      end
      _zz_PerformanceCounterPlugin_logic_branchMissEvent <= (CommitPlugin_logic_commit_reschedulePort_valid && (CommitPlugin_logic_commit_reschedulePort_payload_reason == 8'h10));
      if(PerformanceCounterPlugin_logic_ignoreNextCommit) begin
        if(when_PerformanceCounterPlugin_l65) begin
          PerformanceCounterPlugin_logic_ignoreNextCommit <= 1'b0;
        end
      end
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded <= (_zz_PerformanceCounterPlugin_logic_fsm_counterReaded + 6'h01);
      PerformanceCounterPlugin_logic_commitCount_regNext <= PerformanceCounterPlugin_logic_commitCount;
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2 <= (_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2 + _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2);
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3 <= (_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3 + _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3);
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4 <= (_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4 + _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4);
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5 <= (_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5 + _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5);
      _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6 <= (_zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6 + _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6);
      if(toplevel_EU0_DivPlugin_logic_div_io_cmd_fire) begin
        EU0_DivPlugin_logic_feed_cmdSent <= 1'b1;
      end
      if(when_DivPlugin_l76) begin
        EU0_DivPlugin_logic_feed_cmdSent <= 1'b0;
      end
      if(AguPlugin_setup_port_valid) begin
        AguPlugin_logic_fired <= 1'b1;
      end
      if(when_AguPlugin_l89) begin
        AguPlugin_logic_fired <= 1'b0;
      end
      EnvCallPlugin_logic_flushes_stateReg <= EnvCallPlugin_logic_flushes_stateNext;
      if(integer_RfTranslationPlugin_logic_init_busy) begin
        integer_RfTranslationPlugin_logic_init_counter <= (integer_RfTranslationPlugin_logic_init_counter + 6'h01);
      end
      if(integer_RfAllocationPlugin_logic_init_busy) begin
        integer_RfAllocationPlugin_logic_init_counter <= (integer_RfAllocationPlugin_logic_init_counter + 7'h01);
      end
      BranchContextPlugin_logic_ptr_commited <= BranchContextPlugin_logic_onCommit_commitedNext;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        BranchContextPlugin_logic_ptr_alloc <= BranchContextPlugin_logic_onCommit_commitedNext;
      end
      HistoryPlugin_logic_onCommit_value <= HistoryPlugin_logic_onCommit_valueNext_2;
      HistoryPlugin_logic_onFetch_value <= HistoryPlugin_logic_onFetch_valueNext;
      HistoryPlugin_logic_update_pushes_0_state <= HistoryPlugin_logic_update_pushes_0_stateNext_1;
      if(FetchCachePlugin_setup_historyJump_valid) begin
        HistoryPlugin_logic_update_pushes_0_state <= FetchCachePlugin_setup_historyJump_payload_history;
      end
      HistoryPlugin_logic_update_pushes_2_state <= HistoryPlugin_logic_update_pushes_2_stateNext_2;
      if(DecoderPredictionPlugin_setup_historyPush_flush) begin
        HistoryPlugin_logic_update_pushes_0_state <= HistoryPlugin_logic_update_pushes_2_stateNext_2;
      end
      if(CommitPlugin_logic_reschedule_reschedulePort_valid) begin
        HistoryPlugin_logic_update_pushes_2_state <= HistoryPlugin_logic_update_rescheduleFlush_newHistory;
        HistoryPlugin_logic_update_pushes_0_state <= HistoryPlugin_logic_update_rescheduleFlush_newHistory;
      end
      if(CommitPlugin_logic_reschedule_reschedulePort_valid) begin
        DecoderPredictionPlugin_logic_ras_ptr_push <= DecoderPredictionPlugin_logic_ras_healPush;
        DecoderPredictionPlugin_logic_ras_ptr_pop <= DecoderPredictionPlugin_logic_ras_healPop;
      end
      Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_0_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_0_allocation) begin
        Lsu2Plugin_logic_lq_regs_0_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_0_redoSet) begin
        Lsu2Plugin_logic_lq_regs_0_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_0_delete) begin
        Lsu2Plugin_logic_lq_regs_0_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_0_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338) begin
        Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_0_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_0_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_0_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_0_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_1_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_1_allocation) begin
        Lsu2Plugin_logic_lq_regs_1_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_1_redoSet) begin
        Lsu2Plugin_logic_lq_regs_1_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_1_delete) begin
        Lsu2Plugin_logic_lq_regs_1_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_1_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_1) begin
        Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_1_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_1_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_1_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_1_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_2_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_2_allocation) begin
        Lsu2Plugin_logic_lq_regs_2_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_2_redoSet) begin
        Lsu2Plugin_logic_lq_regs_2_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_2_delete) begin
        Lsu2Plugin_logic_lq_regs_2_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_2_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_2) begin
        Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_2_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_2_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_2_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_2_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_3_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_3_allocation) begin
        Lsu2Plugin_logic_lq_regs_3_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_3_redoSet) begin
        Lsu2Plugin_logic_lq_regs_3_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_3_delete) begin
        Lsu2Plugin_logic_lq_regs_3_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_3_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_3) begin
        Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_3_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_3_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_3_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_3_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_4_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_4_allocation) begin
        Lsu2Plugin_logic_lq_regs_4_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_4_redoSet) begin
        Lsu2Plugin_logic_lq_regs_4_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_4_delete) begin
        Lsu2Plugin_logic_lq_regs_4_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_4_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_4) begin
        Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_4_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_4_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_4_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_4_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_5_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_5_allocation) begin
        Lsu2Plugin_logic_lq_regs_5_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_5_redoSet) begin
        Lsu2Plugin_logic_lq_regs_5_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_5_delete) begin
        Lsu2Plugin_logic_lq_regs_5_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_5_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_5) begin
        Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_5_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_5_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_5_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_5_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_6_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_6_allocation) begin
        Lsu2Plugin_logic_lq_regs_6_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_6_redoSet) begin
        Lsu2Plugin_logic_lq_regs_6_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_6_delete) begin
        Lsu2Plugin_logic_lq_regs_6_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_6_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_6) begin
        Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_6_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_6_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_6_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_6_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_7_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_7_allocation) begin
        Lsu2Plugin_logic_lq_regs_7_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_7_redoSet) begin
        Lsu2Plugin_logic_lq_regs_7_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_7_delete) begin
        Lsu2Plugin_logic_lq_regs_7_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_7_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_7) begin
        Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_7_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_7_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_7_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_7_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_8_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_8_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_8_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_8_allocation) begin
        Lsu2Plugin_logic_lq_regs_8_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_8_redoSet) begin
        Lsu2Plugin_logic_lq_regs_8_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_8_delete) begin
        Lsu2Plugin_logic_lq_regs_8_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_8_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_8) begin
        Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_8_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_8_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_8_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_8_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_9_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_9_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_9_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_9_allocation) begin
        Lsu2Plugin_logic_lq_regs_9_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_9_redoSet) begin
        Lsu2Plugin_logic_lq_regs_9_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_9_delete) begin
        Lsu2Plugin_logic_lq_regs_9_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_9_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_9) begin
        Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_9_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_9_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_9_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_9_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_10_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_10_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_10_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_10_allocation) begin
        Lsu2Plugin_logic_lq_regs_10_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_10_redoSet) begin
        Lsu2Plugin_logic_lq_regs_10_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_10_delete) begin
        Lsu2Plugin_logic_lq_regs_10_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_10_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_10) begin
        Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_10_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_10_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_10_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_10_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_11_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_11_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_11_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_11_allocation) begin
        Lsu2Plugin_logic_lq_regs_11_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_11_redoSet) begin
        Lsu2Plugin_logic_lq_regs_11_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_11_delete) begin
        Lsu2Plugin_logic_lq_regs_11_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_11_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_11) begin
        Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_11_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_11_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_11_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_11_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_12_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_12_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_12_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_12_allocation) begin
        Lsu2Plugin_logic_lq_regs_12_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_12_redoSet) begin
        Lsu2Plugin_logic_lq_regs_12_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_12_delete) begin
        Lsu2Plugin_logic_lq_regs_12_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_12_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_12) begin
        Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_12_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_12_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_12_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_12_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_13_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_13_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_13_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_13_allocation) begin
        Lsu2Plugin_logic_lq_regs_13_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_13_redoSet) begin
        Lsu2Plugin_logic_lq_regs_13_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_13_delete) begin
        Lsu2Plugin_logic_lq_regs_13_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_13_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_13) begin
        Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_13_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_13_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_13_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_13_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_14_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_14_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_14_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_14_allocation) begin
        Lsu2Plugin_logic_lq_regs_14_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_14_redoSet) begin
        Lsu2Plugin_logic_lq_regs_14_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_14_delete) begin
        Lsu2Plugin_logic_lq_regs_14_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_14_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_14) begin
        Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_14_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_14_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_14_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_14_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefill <= (Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefill | Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefillSet);
      Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAny || Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAnySet);
      Lsu2Plugin_logic_lq_regs_15_waitOn_sqWriteback <= (Lsu2Plugin_logic_lq_regs_15_waitOn_sqWriteback || Lsu2Plugin_logic_lq_regs_15_waitOn_sqWritebackSet);
      Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeed <= (Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeed || Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeedSet);
      if(Lsu2Plugin_logic_lq_regs_15_allocation) begin
        Lsu2Plugin_logic_lq_regs_15_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_15_redoSet) begin
        Lsu2Plugin_logic_lq_regs_15_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_lq_regs_15_delete) begin
        Lsu2Plugin_logic_lq_regs_15_valid <= 1'b0;
        Lsu2Plugin_logic_lq_regs_15_redo <= 1'b0;
      end
      if(when_Lsu2Plugin_l338_15) begin
        Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefill <= 2'b00;
        Lsu2Plugin_logic_lq_regs_15_waitOn_cacheRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_15_waitOn_mmuRefillAny <= 1'b0;
        Lsu2Plugin_logic_lq_regs_15_waitOn_sqFeed <= 1'b0;
        Lsu2Plugin_logic_lq_regs_15_waitOn_sqWriteback <= 1'b0;
      end
      Lsu2Plugin_logic_lq_tracker_free <= Lsu2Plugin_logic_lq_tracker_freeNext;
      Lsu2Plugin_logic_lq_ptr_priority <= Lsu2Plugin_logic_lq_onCommit_priority_2;
      Lsu2Plugin_logic_lq_ptr_free <= (Lsu2Plugin_logic_lq_ptr_free + _zz_Lsu2Plugin_logic_lq_ptr_free);
      if(Lsu2Plugin_logic_lq_reservation_kill) begin
        Lsu2Plugin_logic_lq_reservation_valid <= 1'b0;
      end
      if(when_Lsu2Plugin_l484) begin
        Lsu2Plugin_logic_lq_reservation_valid <= 1'b0;
      end else begin
        Lsu2Plugin_logic_lq_reservation_counter <= (Lsu2Plugin_logic_lq_reservation_counter + 7'h01);
      end
      Lsu2Plugin_logic_sq_regs_0_commited <= Lsu2Plugin_logic_sq_regs_0_commitedNext;
      Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_0_allocation) begin
        Lsu2Plugin_logic_sq_regs_0_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_0_redoSet) begin
        Lsu2Plugin_logic_sq_regs_0_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_0_delete) begin
        Lsu2Plugin_logic_sq_regs_0_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_0_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_0_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385) begin
        Lsu2Plugin_logic_sq_regs_0_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_1_commited <= Lsu2Plugin_logic_sq_regs_1_commitedNext;
      Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_1_allocation) begin
        Lsu2Plugin_logic_sq_regs_1_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_1_redoSet) begin
        Lsu2Plugin_logic_sq_regs_1_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_1_delete) begin
        Lsu2Plugin_logic_sq_regs_1_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_1_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_1_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_1) begin
        Lsu2Plugin_logic_sq_regs_1_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_2_commited <= Lsu2Plugin_logic_sq_regs_2_commitedNext;
      Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_2_allocation) begin
        Lsu2Plugin_logic_sq_regs_2_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_2_redoSet) begin
        Lsu2Plugin_logic_sq_regs_2_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_2_delete) begin
        Lsu2Plugin_logic_sq_regs_2_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_2_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_2_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_2) begin
        Lsu2Plugin_logic_sq_regs_2_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_3_commited <= Lsu2Plugin_logic_sq_regs_3_commitedNext;
      Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_3_allocation) begin
        Lsu2Plugin_logic_sq_regs_3_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_3_redoSet) begin
        Lsu2Plugin_logic_sq_regs_3_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_3_delete) begin
        Lsu2Plugin_logic_sq_regs_3_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_3_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_3_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_3) begin
        Lsu2Plugin_logic_sq_regs_3_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_4_commited <= Lsu2Plugin_logic_sq_regs_4_commitedNext;
      Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_4_allocation) begin
        Lsu2Plugin_logic_sq_regs_4_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_4_redoSet) begin
        Lsu2Plugin_logic_sq_regs_4_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_4_delete) begin
        Lsu2Plugin_logic_sq_regs_4_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_4_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_4_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_4) begin
        Lsu2Plugin_logic_sq_regs_4_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_5_commited <= Lsu2Plugin_logic_sq_regs_5_commitedNext;
      Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_5_allocation) begin
        Lsu2Plugin_logic_sq_regs_5_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_5_redoSet) begin
        Lsu2Plugin_logic_sq_regs_5_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_5_delete) begin
        Lsu2Plugin_logic_sq_regs_5_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_5_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_5_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_5) begin
        Lsu2Plugin_logic_sq_regs_5_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_6_commited <= Lsu2Plugin_logic_sq_regs_6_commitedNext;
      Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_6_allocation) begin
        Lsu2Plugin_logic_sq_regs_6_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_6_redoSet) begin
        Lsu2Plugin_logic_sq_regs_6_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_6_delete) begin
        Lsu2Plugin_logic_sq_regs_6_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_6_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_6_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_6) begin
        Lsu2Plugin_logic_sq_regs_6_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_7_commited <= Lsu2Plugin_logic_sq_regs_7_commitedNext;
      Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_7_allocation) begin
        Lsu2Plugin_logic_sq_regs_7_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_7_redoSet) begin
        Lsu2Plugin_logic_sq_regs_7_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_7_delete) begin
        Lsu2Plugin_logic_sq_regs_7_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_7_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_7_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_7) begin
        Lsu2Plugin_logic_sq_regs_7_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_8_commited <= Lsu2Plugin_logic_sq_regs_8_commitedNext;
      Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_8_allocation) begin
        Lsu2Plugin_logic_sq_regs_8_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_8_redoSet) begin
        Lsu2Plugin_logic_sq_regs_8_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_8_delete) begin
        Lsu2Plugin_logic_sq_regs_8_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_8_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_8_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_8) begin
        Lsu2Plugin_logic_sq_regs_8_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_9_commited <= Lsu2Plugin_logic_sq_regs_9_commitedNext;
      Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_9_allocation) begin
        Lsu2Plugin_logic_sq_regs_9_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_9_redoSet) begin
        Lsu2Plugin_logic_sq_regs_9_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_9_delete) begin
        Lsu2Plugin_logic_sq_regs_9_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_9_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_9_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_9) begin
        Lsu2Plugin_logic_sq_regs_9_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_10_commited <= Lsu2Plugin_logic_sq_regs_10_commitedNext;
      Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_10_allocation) begin
        Lsu2Plugin_logic_sq_regs_10_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_10_redoSet) begin
        Lsu2Plugin_logic_sq_regs_10_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_10_delete) begin
        Lsu2Plugin_logic_sq_regs_10_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_10_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_10_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_10) begin
        Lsu2Plugin_logic_sq_regs_10_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_11_commited <= Lsu2Plugin_logic_sq_regs_11_commitedNext;
      Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_11_allocation) begin
        Lsu2Plugin_logic_sq_regs_11_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_11_redoSet) begin
        Lsu2Plugin_logic_sq_regs_11_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_11_delete) begin
        Lsu2Plugin_logic_sq_regs_11_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_11_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_11_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_11) begin
        Lsu2Plugin_logic_sq_regs_11_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_12_commited <= Lsu2Plugin_logic_sq_regs_12_commitedNext;
      Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_12_allocation) begin
        Lsu2Plugin_logic_sq_regs_12_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_12_redoSet) begin
        Lsu2Plugin_logic_sq_regs_12_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_12_delete) begin
        Lsu2Plugin_logic_sq_regs_12_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_12_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_12_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_12) begin
        Lsu2Plugin_logic_sq_regs_12_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_13_commited <= Lsu2Plugin_logic_sq_regs_13_commitedNext;
      Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_13_allocation) begin
        Lsu2Plugin_logic_sq_regs_13_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_13_redoSet) begin
        Lsu2Plugin_logic_sq_regs_13_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_13_delete) begin
        Lsu2Plugin_logic_sq_regs_13_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_13_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_13_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_13) begin
        Lsu2Plugin_logic_sq_regs_13_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_14_commited <= Lsu2Plugin_logic_sq_regs_14_commitedNext;
      Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_14_allocation) begin
        Lsu2Plugin_logic_sq_regs_14_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_14_redoSet) begin
        Lsu2Plugin_logic_sq_regs_14_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_14_delete) begin
        Lsu2Plugin_logic_sq_regs_14_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_14_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_14_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_14) begin
        Lsu2Plugin_logic_sq_regs_14_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_regs_15_commited <= Lsu2Plugin_logic_sq_regs_15_commitedNext;
      Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAny <= (Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAny || Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAnySet);
      if(Lsu2Plugin_logic_sq_regs_15_allocation) begin
        Lsu2Plugin_logic_sq_regs_15_valid <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_15_redoSet) begin
        Lsu2Plugin_logic_sq_regs_15_redo <= 1'b1;
      end
      if(Lsu2Plugin_logic_sq_regs_15_delete) begin
        Lsu2Plugin_logic_sq_regs_15_valid <= 1'b0;
        Lsu2Plugin_logic_sq_regs_15_redo <= 1'b0;
        Lsu2Plugin_logic_sq_regs_15_commited <= 1'b0;
      end
      if(when_Lsu2Plugin_l385_15) begin
        Lsu2Plugin_logic_sq_regs_15_waitOn_mmuRefillAny <= 1'b0;
      end
      Lsu2Plugin_logic_sq_ptr_commit <= Lsu2Plugin_logic_sq_ptr_commitNext;
      Lsu2Plugin_logic_sq_ptr_onFreeLast_valid <= Lsu2Plugin_logic_sq_ptr_onFree_valid;
      Lsu2Plugin_logic_sq_tracker_free <= Lsu2Plugin_logic_sq_tracker_freeNext;
      if(FrontendPlugin_dispatch_isFireing) begin
        Lsu2Plugin_logic_lq_ptr_alloc <= Lsu2Plugin_logic_allocation_loads_alloc_2;
        Lsu2Plugin_logic_sq_ptr_alloc <= Lsu2Plugin_logic_allocation_stores_alloc_2;
      end
      if(Lsu2Plugin_logic_lqSqArbitration_s0_ready) begin
        if(Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT) begin
          if(Lsu2Plugin_logic_lqSqArbitration_s0_LQ_OH[0]) begin
            Lsu2Plugin_logic_lq_regs_0_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID) begin
            Lsu2Plugin_logic_lq_regs_1_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_1) begin
            Lsu2Plugin_logic_lq_regs_2_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_2) begin
            Lsu2Plugin_logic_lq_regs_3_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_3) begin
            Lsu2Plugin_logic_lq_regs_4_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_4) begin
            Lsu2Plugin_logic_lq_regs_5_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_5) begin
            Lsu2Plugin_logic_lq_regs_6_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_6) begin
            Lsu2Plugin_logic_lq_regs_7_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_7) begin
            Lsu2Plugin_logic_lq_regs_8_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_8) begin
            Lsu2Plugin_logic_lq_regs_9_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_9) begin
            Lsu2Plugin_logic_lq_regs_10_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_10) begin
            Lsu2Plugin_logic_lq_regs_11_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_11) begin
            Lsu2Plugin_logic_lq_regs_12_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_12) begin
            Lsu2Plugin_logic_lq_regs_13_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_13) begin
            Lsu2Plugin_logic_lq_regs_14_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID_14) begin
            Lsu2Plugin_logic_lq_regs_15_redo <= 1'b0;
          end
        end
        if(Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT) begin
          if(Lsu2Plugin_logic_lqSqArbitration_s0_SQ_OH[0]) begin
            Lsu2Plugin_logic_sq_regs_0_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID) begin
            Lsu2Plugin_logic_sq_regs_1_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_1) begin
            Lsu2Plugin_logic_sq_regs_2_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_2) begin
            Lsu2Plugin_logic_sq_regs_3_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_3) begin
            Lsu2Plugin_logic_sq_regs_4_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_4) begin
            Lsu2Plugin_logic_sq_regs_5_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_5) begin
            Lsu2Plugin_logic_sq_regs_6_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_6) begin
            Lsu2Plugin_logic_sq_regs_7_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_7) begin
            Lsu2Plugin_logic_sq_regs_8_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_8) begin
            Lsu2Plugin_logic_sq_regs_9_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_9) begin
            Lsu2Plugin_logic_sq_regs_10_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_10) begin
            Lsu2Plugin_logic_sq_regs_11_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_11) begin
            Lsu2Plugin_logic_sq_regs_12_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_12) begin
            Lsu2Plugin_logic_sq_regs_13_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_13) begin
            Lsu2Plugin_logic_sq_regs_14_redo <= 1'b0;
          end
          if(_zz_Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID_14) begin
            Lsu2Plugin_logic_sq_regs_15_redo <= 1'b0;
          end
        end
      end
      if(Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap) begin
        Lsu2Plugin_logic_sharedPip_speculativeHitPredictionGotReschedule <= 1'b0;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_sharedPip_speculativeHitPredictionGotReschedule <= 1'b1;
      end
      if(Lsu2Plugin_logic_sharedPip_hadSpeculativeHitTrap) begin
        Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled <= 1'b0;
      end
      if(Lsu2Plugin_logic_sharedPip_speculateHitTrapRecovered) begin
        Lsu2Plugin_logic_sharedPip_speculativeHitPredictionEnabled <= 1'b1;
      end
      if(when_Lsu2Plugin_l841) begin
        if(when_Lsu2Plugin_l843) begin
          if(Lsu2Plugin_logic_sharedPip_stages_0_feed_TAKE_LQ) begin
            Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask <= 1'b0;
          end
          if(when_Lsu2Plugin_l845) begin
            Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask <= 1'b0;
          end
        end
      end
      if(when_Lsu2Plugin_l849) begin
        Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_lqMask <= 1'b1;
        Lsu2Plugin_logic_sharedPip_feed_lqSqSerializer_sqMask <= 1'b1;
      end
      if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
        case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
          Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
          end
          Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
          end
          Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
          end
          Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          end
          Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
          end
          Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
          end
          Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
          end
          default : begin
            if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
              if(when_Lsu2Plugin_l1333) begin
                if(Lsu2Plugin_logic_sharedPip_stages_3_LR) begin
                  Lsu2Plugin_logic_lq_reservation_valid <= (! Lsu2Plugin_logic_lq_reservation_valid);
                  Lsu2Plugin_logic_lq_reservation_counter <= 7'h00;
                end
              end
            end
          end
        endcase
      end
      Lsu2Plugin_logic_writeback_waitOn_refillSlot <= ((Lsu2Plugin_logic_writeback_waitOn_refillSlot | Lsu2Plugin_logic_writeback_waitOn_refillSlotSet) & (~ DataCachePlugin_setup_refillCompletions));
      Lsu2Plugin_logic_writeback_waitOn_refillSlotAny <= ((Lsu2Plugin_logic_writeback_waitOn_refillSlotAny || Lsu2Plugin_logic_writeback_waitOn_refillSlotAnySet) && (! (|DataCachePlugin_setup_refillCompletions)));
      if(Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready) begin
        toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rValid <= Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_valid;
      end
      Lsu2Plugin_logic_sq_ptr_writeBack <= (Lsu2Plugin_logic_sq_ptr_writeBack + _zz_Lsu2Plugin_logic_sq_ptr_writeBack);
      Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_valid <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_valid;
      if(when_Lsu2Plugin_l1488) begin
        if(Lsu2Plugin_logic_writeback_rsp_delayed_1_payload_redo) begin
          Lsu2Plugin_logic_writeback_generation <= (! Lsu2Plugin_logic_writeback_generation);
          Lsu2Plugin_logic_sq_ptr_writeBack <= Lsu2Plugin_logic_sq_ptr_free;
        end
      end
      if(when_Lsu2Plugin_l1509) begin
        Lsu2Plugin_logic_sq_ptr_writeBack <= (Lsu2Plugin_logic_sq_ptr_writeBack + 5'h01);
      end
      if(Lsu2Plugin_logic_sq_ptr_onFree_valid) begin
        Lsu2Plugin_logic_sq_ptr_free <= (Lsu2Plugin_logic_sq_ptr_free + 5'h01);
        Lsu2Plugin_logic_sq_ptr_priority <= (Lsu2Plugin_logic_sq_ptr_priority <<< 1);
        if(when_Lsu2Plugin_l1521) begin
          Lsu2Plugin_logic_sq_ptr_priority <= 15'h7fff;
        end
      end
      Lsu2Plugin_logic_flush_doit <= (Lsu2Plugin_logic_sq_ptr_commit == Lsu2Plugin_logic_sq_ptr_free);
      if(Lsu2Plugin_setup_flushPort_cmd_valid) begin
        Lsu2Plugin_logic_flush_busy <= 1'b1;
        Lsu2Plugin_logic_flush_doit <= 1'b0;
      end
      if(when_Lsu2Plugin_l1553) begin
        if(when_Lsu2Plugin_l1561) begin
          if(Lsu2Plugin_setup_cacheStore_rsp_payload_redo) begin
            Lsu2Plugin_logic_writeback_generation <= (! Lsu2Plugin_logic_writeback_generation);
          end
        end
        if(when_Lsu2Plugin_l1569) begin
          Lsu2Plugin_logic_flush_busy <= 1'b0;
        end
      end
      LsuPlugin_peripheralBus_rsp_valid_regNext <= LsuPlugin_peripheralBus_rsp_valid;
      if(Lsu2Plugin_logic_special_hit) begin
        Lsu2Plugin_logic_special_enabled <= 1'b1;
      end
      if(Lsu2Plugin_logic_special_fire) begin
        Lsu2Plugin_logic_special_enabled <= 1'b0;
      end
      if(LsuPlugin_peripheralBus_cmd_fire) begin
        Lsu2Plugin_logic_special_cmdSent <= 1'b1;
      end
      if(Lsu2Plugin_logic_special_fire) begin
        Lsu2Plugin_logic_special_cmdSent <= 1'b0;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_lq_ptr_free <= 5'h00;
        Lsu2Plugin_logic_lq_ptr_alloc <= 5'h00;
        Lsu2Plugin_logic_lq_ptr_priority <= 15'h0000;
        Lsu2Plugin_logic_sq_ptr_alloc <= Lsu2Plugin_logic_sq_ptr_commitNext;
        Lsu2Plugin_logic_special_enabled <= 1'b0;
      end
      if(PrivilegedPlugin_setup_xretAwayFromMachine) begin
        MmuPlugin_logic_status_mprv <= 1'b0;
      end
      FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_value <= FetchCachePlugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
      FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_value <= FetchCachePlugin_setup_translationStorage_logic_sl_1_allocId_valueNext;
      Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_value <= Lsu2Plugin_setup_translationStorage_logic_sl_0_allocId_valueNext;
      Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_value <= Lsu2Plugin_setup_translationStorage_logic_sl_1_allocId_valueNext;
      Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg <= Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL_overloaded;
      if(when_MmuPlugin_l260) begin
        Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_0_reg <= 1'b1;
      end
      Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg <= Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded;
      if(when_MmuPlugin_l260_1) begin
        Lsu2Plugin_logic_sharedPip_translationPort_logic_allowRefillBypass_1_reg <= 1'b1;
      end
      PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt <= PrivilegedPlugin_logic_interrupt_valid;
      if(PrivilegedPlugin_logic_decoderInterrupt_pendingInterrupt) begin
        PrivilegedPlugin_logic_decoderInterrupt_counter <= (PrivilegedPlugin_logic_decoderInterrupt_counter + 3'b001);
      end
      if(when_PrivilegedPlugin_l668) begin
        PrivilegedPlugin_logic_decoderInterrupt_counter <= 3'b000;
      end
      if(when_PrivilegedPlugin_l672) begin
        PrivilegedPlugin_logic_decoderInterrupt_raised <= 1'b1;
      end
      if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_fire) begin
        PerformanceCounterPlugin_logic_csrRead_fired <= 1'b1;
      end
      if(EU0_CsrAccessPlugin_setup_onReadMovingOff) begin
        PerformanceCounterPlugin_logic_csrRead_fired <= 1'b0;
      end
      if(PerformanceCounterPlugin_logic_fsm_csrWriteCmd_fire) begin
        PerformanceCounterPlugin_logic_csrWrite_fired <= 1'b1;
      end
      if(EU0_CsrAccessPlugin_setup_onWriteMovingOff) begin
        PerformanceCounterPlugin_logic_csrWrite_fired <= 1'b0;
      end
      FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg <= FetchPlugin_stages_1_MmuPlugin_logic_ALLOW_REFILL_overloaded;
      if(when_MmuPlugin_l260_2) begin
        FetchCachePlugin_logic_translationPort_logic_allowRefillBypass_0_reg <= 1'b1;
      end
      MmuPlugin_logic_refill_cacheRefill <= ((MmuPlugin_logic_refill_cacheRefill | MmuPlugin_logic_refill_cacheRefillSet) & (~ DataCachePlugin_setup_refillCompletions));
      MmuPlugin_logic_refill_cacheRefillAny <= ((MmuPlugin_logic_refill_cacheRefillAny || MmuPlugin_logic_refill_cacheRefillAnySet) && (! (|DataCachePlugin_setup_refillCompletions)));
      MmuPlugin_logic_refill_load_rsp_valid <= MmuPlugin_setup_cacheLoad_rsp_valid;
      if(MmuPlugin_setup_invalidatePort_cmd_valid) begin
        MmuPlugin_logic_invalidate_requested <= 1'b1;
      end
      if(when_MmuPlugin_l492) begin
        MmuPlugin_logic_invalidate_counter <= (MmuPlugin_logic_invalidate_counter + 6'h01);
      end
      if(when_MmuPlugin_l505) begin
        MmuPlugin_logic_invalidate_counter <= 6'h00;
        MmuPlugin_logic_invalidate_requested <= 1'b0;
      end
      MmuPlugin_logic_invalidate_done_regNext <= MmuPlugin_logic_invalidate_done;
      Lsu2Plugin_logic_sharedPip_stages_1_valid <= _zz_Lsu2Plugin_logic_sharedPip_stages_1_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_sharedPip_stages_1_valid <= 1'b0;
      end
      Lsu2Plugin_logic_sharedPip_stages_2_valid <= Lsu2Plugin_logic_sharedPip_stages_1_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_sharedPip_stages_2_valid <= 1'b0;
      end
      Lsu2Plugin_logic_sharedPip_stages_3_valid <= Lsu2Plugin_logic_sharedPip_stages_2_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_sharedPip_stages_3_valid <= 1'b0;
      end
      if(Lsu2Plugin_logic_lqSqArbitration_s0_ready_output) begin
        Lsu2Plugin_logic_lqSqArbitration_s1_valid <= Lsu2Plugin_logic_lqSqArbitration_s0_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        Lsu2Plugin_logic_lqSqArbitration_s1_valid <= 1'b0;
      end
      Lsu2Plugin_logic_special_atomic_stateReg <= Lsu2Plugin_logic_special_atomic_stateNext;
      (* parallel_case *)
      case(1) // synthesis parallel_case
        (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
        end
        (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
        end
        (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
          if(Lsu2Plugin_setup_cacheLoad_rsp_valid) begin
            Lsu2Plugin_logic_special_atomic_comp_rfWrite <= 1'b0;
          end
        end
        (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
          Lsu2Plugin_logic_special_atomic_lockDelayCounter <= (Lsu2Plugin_logic_special_atomic_lockDelayCounter + 2'b01);
        end
        (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
        end
        (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
          Lsu2Plugin_logic_special_atomic_comp_wakeRf <= 1'b0;
          Lsu2Plugin_logic_special_atomic_comp_rfWrite <= 1'b0;
        end
        (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
        end
        (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l253) begin
        Lsu2Plugin_logic_special_atomic_comp_rfWrite <= Lsu2Plugin_logic_sq_mem_writeRd;
      end
      if(when_StateMachine_l253_1) begin
        Lsu2Plugin_logic_special_atomic_comp_wakeRf <= Lsu2Plugin_logic_sq_mem_writeRd;
        Lsu2Plugin_logic_special_atomic_comp_rfWrite <= (Lsu2Plugin_logic_special_storeSc && Lsu2Plugin_logic_sq_mem_writeRd);
      end
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_stateNext;
      if(when_CsrRamPlugin_l61) begin
        CsrRamPlugin_logic_flush_counter <= (CsrRamPlugin_logic_flush_counter + 6'h01);
      end
      if(when_CsrAccessPlugin_l326) begin
        PrivilegedPlugin_logic_machine_cause_interrupt <= EU0_CsrAccessPlugin_setup_onWriteBits[31];
        PrivilegedPlugin_logic_machine_cause_code <= EU0_CsrAccessPlugin_setup_onWriteBits[3 : 0];
      end
      if(when_CsrAccessPlugin_l326_1) begin
        PrivilegedPlugin_logic_machine_mstatus_mpp <= EU0_CsrAccessPlugin_setup_onWriteBits[12 : 11];
        PrivilegedPlugin_logic_machine_mstatus_mpie <= EU0_CsrAccessPlugin_setup_onWriteBits[7];
        PrivilegedPlugin_logic_machine_mstatus_mie <= EU0_CsrAccessPlugin_setup_onWriteBits[3];
        PrivilegedPlugin_logic_machine_mstatus_fs <= EU0_CsrAccessPlugin_setup_onWriteBits[14 : 13];
        PrivilegedPlugin_logic_supervisor_sstatus_spp <= EU0_CsrAccessPlugin_setup_onWriteBits[8 : 8];
        PrivilegedPlugin_logic_supervisor_sstatus_spie <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_supervisor_sstatus_sie <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
        MmuPlugin_logic_status_mxr <= EU0_CsrAccessPlugin_setup_onWriteBits[19];
        MmuPlugin_logic_status_sum <= EU0_CsrAccessPlugin_setup_onWriteBits[18];
        MmuPlugin_logic_status_mprv <= EU0_CsrAccessPlugin_setup_onWriteBits[17];
      end
      if(when_CsrAccessPlugin_l326_2) begin
        PrivilegedPlugin_logic_supervisor_sip_seipSoft <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        PrivilegedPlugin_logic_supervisor_sip_stip <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_supervisor_sip_ssip <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
      end
      if(when_CsrAccessPlugin_l326_3) begin
        PrivilegedPlugin_logic_machine_mie_meie <= EU0_CsrAccessPlugin_setup_onWriteBits[11];
        PrivilegedPlugin_logic_machine_mie_mtie <= EU0_CsrAccessPlugin_setup_onWriteBits[7];
        PrivilegedPlugin_logic_machine_mie_msie <= EU0_CsrAccessPlugin_setup_onWriteBits[3];
        PrivilegedPlugin_logic_supervisor_sie_seie <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        PrivilegedPlugin_logic_supervisor_sie_stie <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_supervisor_sie_ssie <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
      end
      if(when_CsrAccessPlugin_l326_4) begin
        PrivilegedPlugin_logic_machine_medeleg_iam <= EU0_CsrAccessPlugin_setup_onWriteBits[0];
        PrivilegedPlugin_logic_machine_medeleg_bp <= EU0_CsrAccessPlugin_setup_onWriteBits[3];
        PrivilegedPlugin_logic_machine_medeleg_eu <= EU0_CsrAccessPlugin_setup_onWriteBits[8];
        PrivilegedPlugin_logic_machine_medeleg_es <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        PrivilegedPlugin_logic_machine_medeleg_ipf <= EU0_CsrAccessPlugin_setup_onWriteBits[12];
        PrivilegedPlugin_logic_machine_medeleg_lpf <= EU0_CsrAccessPlugin_setup_onWriteBits[13];
        PrivilegedPlugin_logic_machine_medeleg_spf <= EU0_CsrAccessPlugin_setup_onWriteBits[15];
      end
      if(when_CsrAccessPlugin_l326_5) begin
        PrivilegedPlugin_logic_machine_mideleg_se <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        PrivilegedPlugin_logic_machine_mideleg_st <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_machine_mideleg_ss <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
      end
      if(when_CsrAccessPlugin_l326_6) begin
        PrivilegedPlugin_logic_supervisor_cause_interrupt <= EU0_CsrAccessPlugin_setup_onWriteBits[31];
        PrivilegedPlugin_logic_supervisor_cause_code <= EU0_CsrAccessPlugin_setup_onWriteBits[3 : 0];
      end
      if(when_CsrAccessPlugin_l326_7) begin
        PrivilegedPlugin_logic_supervisor_sstatus_spp <= EU0_CsrAccessPlugin_setup_onWriteBits[8 : 8];
        PrivilegedPlugin_logic_supervisor_sstatus_spie <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        PrivilegedPlugin_logic_supervisor_sstatus_sie <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
        PrivilegedPlugin_logic_machine_mstatus_fs <= EU0_CsrAccessPlugin_setup_onWriteBits[14 : 13];
        MmuPlugin_logic_status_mxr <= EU0_CsrAccessPlugin_setup_onWriteBits[19];
        MmuPlugin_logic_status_sum <= EU0_CsrAccessPlugin_setup_onWriteBits[18];
      end
      if(when_CsrAccessPlugin_l326_8) begin
        if(PrivilegedPlugin_logic_machine_mideleg_se) begin
          PrivilegedPlugin_logic_supervisor_sie_seie <= EU0_CsrAccessPlugin_setup_onWriteBits[9];
        end
        if(PrivilegedPlugin_logic_machine_mideleg_st) begin
          PrivilegedPlugin_logic_supervisor_sie_stie <= EU0_CsrAccessPlugin_setup_onWriteBits[5];
        end
        if(PrivilegedPlugin_logic_machine_mideleg_ss) begin
          PrivilegedPlugin_logic_supervisor_sie_ssie <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
        end
      end
      if(when_CsrAccessPlugin_l326_9) begin
        if(PrivilegedPlugin_logic_machine_mideleg_ss) begin
          PrivilegedPlugin_logic_supervisor_sip_ssip <= EU0_CsrAccessPlugin_setup_onWriteBits[1];
        end
      end
      if(when_CsrAccessPlugin_l326_10) begin
        _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_7 <= EU0_CsrAccessPlugin_setup_onWriteBits[2 : 0];
      end
      if(when_CsrAccessPlugin_l326_11) begin
        _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_8 <= EU0_CsrAccessPlugin_setup_onWriteBits[2 : 0];
      end
      if(when_CsrAccessPlugin_l326_12) begin
        _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_9 <= EU0_CsrAccessPlugin_setup_onWriteBits[2 : 0];
      end
      if(when_CsrAccessPlugin_l326_13) begin
        _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_10 <= EU0_CsrAccessPlugin_setup_onWriteBits[2 : 0];
      end
      if(when_CsrAccessPlugin_l331) begin
        if(when_CsrAccessPlugin_l326_14) begin
          MmuPlugin_logic_satp_mode <= EU0_CsrAccessPlugin_setup_onWriteBits[31 : 31];
          MmuPlugin_logic_satp_ppn <= EU0_CsrAccessPlugin_setup_onWriteBits[19 : 0];
        end
      end
      if(when_CsrAccessPlugin_l336) begin
        EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired <= 1'b1;
      end
      if(EU0_CsrAccessPlugin_setup_onWriteMovingOff) begin
        EU0_CsrAccessPlugin_logic_fsm_writeLogic_ramWrite_fired <= 1'b0;
      end
      EU0_CsrAccessPlugin_logic_fsm_stateReg <= EU0_CsrAccessPlugin_logic_fsm_stateNext;
      if(DecoderPlugin_logic_exception_set) begin
        DecoderPlugin_logic_exception_trigged <= 1'b1;
      end
      if(DecoderPlugin_logic_exception_clear) begin
        DecoderPlugin_logic_exception_trigged <= 1'b0;
      end
      DecoderPlugin_logic_exception_doItAgain <= DecoderPlugin_logic_exception_doIt;
      FrontendPlugin_decoded_OP_ID <= (FrontendPlugin_decoded_OP_ID + _zz_FrontendPlugin_decoded_OP_ID);
      if(FrontendPlugin_serialized_valid) begin
        DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle <= 1'b0;
      end
      if(when_DecoderPredictionPlugin_l236) begin
        DecoderPredictionPlugin_logic_decodePatch_applyIt_firstCycle <= 1'b1;
      end
      ALU0_ExecutionUnitBase_pipeline_fetch_1_valid <= ALU0_ExecutionUnitBase_pipeline_fetch_0_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        ALU0_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      end
      ALU0_ExecutionUnitBase_pipeline_execute_1_valid <= ALU0_ExecutionUnitBase_pipeline_execute_0_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        ALU0_ExecutionUnitBase_pipeline_execute_1_valid <= 1'b0;
      end
      ALU1_ExecutionUnitBase_pipeline_fetch_1_valid <= ALU1_ExecutionUnitBase_pipeline_fetch_0_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        ALU1_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      end
      ALU1_ExecutionUnitBase_pipeline_execute_1_valid <= ALU1_ExecutionUnitBase_pipeline_execute_0_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        ALU1_ExecutionUnitBase_pipeline_execute_1_valid <= 1'b0;
      end
      if(EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output) begin
        EU0_ExecutionUnitBase_pipeline_fetch_1_valid <= EU0_ExecutionUnitBase_pipeline_fetch_0_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        EU0_ExecutionUnitBase_pipeline_fetch_1_valid <= 1'b0;
      end
      if(EU0_ExecutionUnitBase_pipeline_execute_0_ready_output) begin
        EU0_ExecutionUnitBase_pipeline_execute_1_valid <= _zz_EU0_ExecutionUnitBase_pipeline_execute_1_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        EU0_ExecutionUnitBase_pipeline_execute_1_valid <= 1'b0;
      end
      if(EU0_ExecutionUnitBase_pipeline_execute_1_ready_output) begin
        EU0_ExecutionUnitBase_pipeline_execute_2_valid <= _zz_EU0_ExecutionUnitBase_pipeline_execute_2_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        EU0_ExecutionUnitBase_pipeline_execute_2_valid <= 1'b0;
      end
      if(BranchContextPlugin_free_learn_valid) begin
        BranchContextPlugin_logic_ptr_free <= (BranchContextPlugin_logic_ptr_free + 5'h01);
      end
      if(toplevel_DispatchPlugin_logic_queue_io_push_fire) begin
        DispatchPlugin_logic_ptr_next <= (DispatchPlugin_logic_ptr_next + 6'h02);
        DispatchPlugin_logic_ptr_current <= (DispatchPlugin_logic_ptr_current + 6'h02);
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        DispatchPlugin_logic_ptr_next <= (_zz_DispatchPlugin_logic_ptr_next + 6'h02);
        DispatchPlugin_logic_ptr_current <= (CommitPlugin_logic_commit_reschedulePort_payload_robIdNext - 6'h20);
      end
      if(when_DispatchPlugin_l192) begin
        DispatchPlugin_logic_push_fenceYoungerLast <= DispatchPlugin_logic_push_fenceYounger;
      end
      DispatchPlugin_logic_pop_0_stagesList_1_valid <= DispatchPlugin_logic_pop_0_stagesList_0_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        DispatchPlugin_logic_pop_0_stagesList_1_valid <= 1'b0;
      end
      DispatchPlugin_logic_pop_1_stagesList_1_valid <= DispatchPlugin_logic_pop_1_stagesList_0_valid;
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        DispatchPlugin_logic_pop_1_stagesList_1_valid <= 1'b0;
      end
      if(DispatchPlugin_logic_pop_2_stagesList_0_ready_output) begin
        DispatchPlugin_logic_pop_2_stagesList_1_valid <= DispatchPlugin_logic_pop_2_stagesList_0_valid;
      end
      if(CommitPlugin_logic_commit_reschedulePort_valid) begin
        DispatchPlugin_logic_pop_2_stagesList_1_valid <= 1'b0;
      end
      if(RfDependencyPlugin_logic_forRf_integer_init_busy) begin
        RfDependencyPlugin_logic_forRf_integer_init_counter <= (RfDependencyPlugin_logic_forRf_integer_init_counter + 7'h01);
      end
      if(FrontendPlugin_allocated_ready_output) begin
        FrontendPlugin_dispatch_valid <= _zz_FrontendPlugin_dispatch_valid;
      end
      if(CommitPlugin_logic_reschedule_reschedulePort_valid) begin
        FrontendPlugin_dispatch_valid <= 1'b0;
      end
      if(FrontendPlugin_decoded_ready_output) begin
        FrontendPlugin_serialized_valid <= _zz_FrontendPlugin_serialized_valid;
      end
      if(when_Connection_l66) begin
        FrontendPlugin_serialized_valid <= 1'b0;
      end
      PcPlugin_logic_init_counter <= (PcPlugin_logic_init_counter + _zz_PcPlugin_logic_init_counter);
      if(PcPlugin_logic_fetchPc_correction) begin
        PcPlugin_logic_fetchPc_correctionReg <= 1'b1;
      end
      if(PcPlugin_logic_fetchPc_output_fire) begin
        PcPlugin_logic_fetchPc_correctionReg <= 1'b0;
      end
      if(when_PcPlugin_l82) begin
        PcPlugin_logic_fetchPc_inc <= 1'b0;
      end
      if(PcPlugin_logic_fetchPc_output_fire) begin
        PcPlugin_logic_fetchPc_inc <= 1'b1;
      end
      if(when_PcPlugin_l82_1) begin
        PcPlugin_logic_fetchPc_inc <= 1'b0;
      end
      if(when_PcPlugin_l98) begin
        PcPlugin_logic_fetchPc_pcReg <= PcPlugin_logic_fetchPc_pc;
      end
      if(when_Connection_l54) begin
        FetchPlugin_stages_1_valid <= 1'b0;
      end
      if(FetchPlugin_stages_0_ready_output) begin
        FetchPlugin_stages_1_valid <= _zz_FetchPlugin_stages_1_valid;
      end
      if(FetchPlugin_stages_1_ready_output) begin
        FetchPlugin_stages_2_valid <= _zz_FetchPlugin_stages_2_valid;
      end
      if(when_Connection_l66_1) begin
        FetchPlugin_stages_2_valid <= 1'b0;
      end
      if(_zz_AlignerPlugin_setup_s2m_valid) begin
        FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid <= 1'b1;
      end
      if(AlignerPlugin_setup_s2m_ready) begin
        FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid <= 1'b0;
      end
      if(FrontendPlugin_aligned_isFlushed) begin
        FetchPlugin_stages_2_to_AlignerPlugin_setup_s2m_rValid <= 1'b0;
      end
      PerformanceCounterPlugin_logic_fsm_stateReg <= PerformanceCounterPlugin_logic_fsm_stateNext;
      case(PerformanceCounterPlugin_logic_fsm_stateReg)
        PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
          if(!PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
            if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
              PerformanceCounterPlugin_logic_fsm_done <= 1'b0;
            end
          end
        end
        PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
        end
        PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
          if(when_PerformanceCounterPlugin_l201) begin
            case(PerformanceCounterPlugin_logic_fsm_cmd_address)
              3'b000 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded[5] <= 1'b0;
              end
              3'b010 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2[5] <= 1'b0;
              end
              3'b011 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3[5] <= 1'b0;
              end
              3'b100 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4[5] <= 1'b0;
              end
              3'b101 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5[5] <= 1'b0;
              end
              3'b110 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6[5] <= 1'b0;
              end
              default : begin
              end
            endcase
          end
          if(!PerformanceCounterPlugin_logic_fsm_cmd_flusher) begin
            PerformanceCounterPlugin_logic_fsm_done <= 1'b1;
          end
        end
        PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
        end
        PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
        end
        PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
        end
        PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
          if(when_PerformanceCounterPlugin_l161) begin
            case(PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address)
              3'b000 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded <= _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded[5:0];
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded[5] <= 1'b0;
              end
              3'b010 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2 <= _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2_1[5:0];
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_2[5] <= 1'b0;
              end
              3'b011 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3 <= _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3_2[5:0];
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_3[5] <= 1'b0;
              end
              3'b100 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4 <= _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4_2[5:0];
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_4[5] <= 1'b0;
              end
              3'b101 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5 <= _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5_2[5:0];
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_5[5] <= 1'b0;
              end
              3'b110 : begin
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6 <= _zz__zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6_2[5:0];
                _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_6[5] <= 1'b0;
              end
              default : begin
              end
            endcase
          end
          if(when_PerformanceCounterPlugin_l169) begin
            PerformanceCounterPlugin_logic_ignoreNextCommit <= 1'b1;
          end
        end
        PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
        end
        default : begin
        end
      endcase
      PrivilegedPlugin_logic_fsm_stateReg <= PrivilegedPlugin_logic_fsm_stateNext;
      case(PrivilegedPlugin_logic_fsm_stateReg)
        PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
          PrivilegedPlugin_setup_privilege <= PrivilegedPlugin_logic_fsm_xret_targetPrivilege;
          case(switch_PrivilegedPlugin_l953)
            2'b11 : begin
              PrivilegedPlugin_logic_machine_mstatus_mpp <= 2'b00;
              PrivilegedPlugin_logic_machine_mstatus_mie <= PrivilegedPlugin_logic_machine_mstatus_mpie;
              PrivilegedPlugin_logic_machine_mstatus_mpie <= 1'b1;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_supervisor_sstatus_spp <= 1'b0;
              PrivilegedPlugin_logic_supervisor_sstatus_sie <= PrivilegedPlugin_logic_supervisor_sstatus_spie;
              PrivilegedPlugin_logic_supervisor_sstatus_spie <= 1'b1;
            end
            default : begin
            end
          endcase
        end
        PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
        end
        PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
          PrivilegedPlugin_setup_privilege <= PrivilegedPlugin_logic_fsm_trap_targetPrivilege;
          case(PrivilegedPlugin_logic_fsm_trap_targetPrivilege)
            2'b11 : begin
              PrivilegedPlugin_logic_machine_mstatus_mie <= 1'b0;
              PrivilegedPlugin_logic_machine_mstatus_mpie <= PrivilegedPlugin_logic_machine_mstatus_mie;
              PrivilegedPlugin_logic_machine_mstatus_mpp <= PrivilegedPlugin_setup_privilege;
              PrivilegedPlugin_logic_machine_cause_interrupt <= PrivilegedPlugin_logic_fsm_trap_interrupt;
              PrivilegedPlugin_logic_machine_cause_code <= PrivilegedPlugin_logic_fsm_trap_code;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_supervisor_sstatus_sie <= 1'b0;
              PrivilegedPlugin_logic_supervisor_sstatus_spie <= PrivilegedPlugin_logic_supervisor_sstatus_sie;
              PrivilegedPlugin_logic_supervisor_sstatus_spp <= PrivilegedPlugin_setup_privilege[0 : 0];
              PrivilegedPlugin_logic_supervisor_cause_interrupt <= PrivilegedPlugin_logic_fsm_trap_interrupt;
              PrivilegedPlugin_logic_supervisor_cause_code <= PrivilegedPlugin_logic_fsm_trap_code;
            end
            default : begin
            end
          endcase
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l253_2) begin
        PrivilegedPlugin_logic_decoderInterrupt_raised <= 1'b0;
      end
      if(FetchCachePlugin_logic_banks_0_read_cmd_valid) begin
        when_MultiportRam_l328 <= (_zz_when_MultiportRam_l328_4 && (FetchCachePlugin_logic_banks_0_write_payload_address == FetchCachePlugin_logic_banks_0_read_cmd_payload));
      end
      if(FetchCachePlugin_logic_banks_1_read_cmd_valid) begin
        when_MultiportRam_l328_1 <= (_zz_when_MultiportRam_l328_3 && (FetchCachePlugin_logic_banks_1_write_payload_address == FetchCachePlugin_logic_banks_1_read_cmd_payload));
      end
      if(FetchCachePlugin_logic_banks_2_read_cmd_valid) begin
        when_MultiportRam_l328_2 <= (_zz_when_MultiportRam_l328_2 && (FetchCachePlugin_logic_banks_2_write_payload_address == FetchCachePlugin_logic_banks_2_read_cmd_payload));
      end
      if(FetchCachePlugin_logic_banks_3_read_cmd_valid) begin
        when_MultiportRam_l328_3 <= (_zz_when_MultiportRam_l328_1 && (FetchCachePlugin_logic_banks_3_write_payload_address == FetchCachePlugin_logic_banks_3_read_cmd_payload));
      end
      if(FetchPlugin_stages_0_ready) begin
        when_MultiportRam_l328_4 <= (_zz_when_MultiportRam_l328 && (GSharePlugin_logic_mem_write_payload_address == FetchPlugin_stages_0_GSharePlugin_logic_HASH));
      end
      if(Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_valid) begin
        when_MultiportRam_l362 <= (_zz_when_MultiportRam_l362_1 && (_zz_when_MultiportRam_l362_2 == Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_payload));
      end
      if(Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_valid) begin
        when_MultiportRam_l362_1 <= (_zz_when_MultiportRam_l362 && (_zz_when_MultiportRam_l362_3 == Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_payload));
      end
    end
  end

  always @(posedge clk) begin
    if(when_FetchCachePlugin_l422) begin
      FetchCachePlugin_logic_refill_address <= FetchCachePlugin_logic_refill_start_address;
      FetchCachePlugin_logic_refill_isIo <= FetchCachePlugin_logic_refill_start_isIo;
      FetchCachePlugin_logic_refill_wayToAllocate <= FetchCachePlugin_logic_refill_start_wayToAllocate;
    end
    if(AlignerPlugin_logic_fireInput) begin
      AlignerPlugin_logic_buffer_data <= AlignerPlugin_setup_s2m_Fetch_WORD;
      AlignerPlugin_logic_buffer_pc <= AlignerPlugin_setup_s2m_Fetch_FETCH_PC;
      AlignerPlugin_logic_buffer_fault <= AlignerPlugin_setup_s2m_Fetch_WORD_FAULT;
      AlignerPlugin_logic_buffer_fault_page <= AlignerPlugin_setup_s2m_Fetch_WORD_FAULT_PAGE;
      AlignerPlugin_logic_buffer_branchValid <= (AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_VALID && (! _zz_FrontendPlugin_aligned_Prediction_ALIGNED_BRANCH_VALID_1));
      AlignerPlugin_logic_buffer_branchSlice <= AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_SLICE;
      AlignerPlugin_logic_buffer_branchPcNext <= AlignerPlugin_setup_s2m_Prediction_WORD_BRANCH_PC_NEXT;
      AlignerPlugin_logic_buffer_wordContexts_0 <= AlignerPlugin_setup_s2m_BRANCH_HISTORY;
      AlignerPlugin_logic_buffer_wordContexts_1 <= AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALID;
      AlignerPlugin_logic_buffer_wordContexts_2 <= AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_SLICE;
      AlignerPlugin_logic_buffer_wordContexts_3 <= AlignerPlugin_setup_s2m_Prediction_BRANCH_HISTORY_PUSH_VALUE;
      AlignerPlugin_logic_buffer_wordContexts_4_0 <= AlignerPlugin_setup_s2m_GSHARE_COUNTER_0;
      AlignerPlugin_logic_buffer_wordContexts_4_1 <= AlignerPlugin_setup_s2m_GSHARE_COUNTER_1;
      AlignerPlugin_logic_buffer_firstWordContexts_0 <= AlignerPlugin_setup_s2m_FETCH_ID;
    end
    CommitPlugin_logic_ptr_robLineMaskRsp <= CommitPlugin_setup_robLineMask_mask;
    if(when_CommitPlugin_l131) begin
      CommitPlugin_logic_reschedule_robId <= ((((_zz_CommitPlugin_logic_reschedule_trap ? _zz_CommitPlugin_logic_reschedule_robId : _zz_CommitPlugin_logic_reschedule_robId_1) | (_zz_CommitPlugin_logic_reschedule_trap_1 ? _zz_CommitPlugin_logic_reschedule_robId_2 : _zz_CommitPlugin_logic_reschedule_robId_3)) | ((_zz_CommitPlugin_logic_reschedule_trap_2 ? _zz_CommitPlugin_logic_reschedule_robId_4 : _zz_CommitPlugin_logic_reschedule_robId_5) | (_zz_CommitPlugin_logic_reschedule_trap_3 ? _zz_CommitPlugin_logic_reschedule_robId_6 : _zz_CommitPlugin_logic_reschedule_robId_7))) | ((_zz_CommitPlugin_logic_reschedule_trap_4 ? EU0_CsrAccessPlugin_setup_trap_payload_robId : 6'h00) | (_zz_CommitPlugin_logic_reschedule_trap_5 ? ALU1_BranchPlugin_setup_reschedule_payload_robId : 6'h00)));
      CommitPlugin_logic_reschedule_trap <= _zz_CommitPlugin_logic_reschedule_trap_6[0];
      CommitPlugin_logic_reschedule_pcTarget <= (((CommitPlugin_logic_reschedule_portsLogic_hits[0] ? Lsu2Plugin_setup_sharedTrap_payload_pcTarget : 32'h00000000) | (CommitPlugin_logic_reschedule_portsLogic_hits[2] ? ALU0_BranchPlugin_setup_reschedule_payload_pcTarget : 32'h00000000)) | (CommitPlugin_logic_reschedule_portsLogic_hits[5] ? ALU1_BranchPlugin_setup_reschedule_payload_pcTarget : 32'h00000000));
      CommitPlugin_logic_reschedule_cause <= ((((_zz_CommitPlugin_logic_reschedule_cause ? _zz_CommitPlugin_logic_reschedule_cause_1 : _zz_CommitPlugin_logic_reschedule_cause_2) | (_zz_CommitPlugin_logic_reschedule_cause_3 ? _zz_CommitPlugin_logic_reschedule_cause_4 : _zz_CommitPlugin_logic_reschedule_cause_5)) | ((_zz_CommitPlugin_logic_reschedule_cause_6 ? _zz_CommitPlugin_logic_reschedule_cause_7 : _zz_CommitPlugin_logic_reschedule_cause_8) | (_zz_CommitPlugin_logic_reschedule_cause_9 ? _zz_CommitPlugin_logic_reschedule_cause_10 : _zz_CommitPlugin_logic_reschedule_cause_11))) | ((CommitPlugin_logic_reschedule_portsLogic_hits[4] ? EU0_CsrAccessPlugin_setup_trap_payload_cause : 4'b0000) | (CommitPlugin_logic_reschedule_portsLogic_hits[5] ? ALU1_BranchPlugin_setup_reschedule_payload_cause : 4'b0000)));
      CommitPlugin_logic_reschedule_reason <= ((((_zz_CommitPlugin_logic_reschedule_reason ? _zz_CommitPlugin_logic_reschedule_reason_1 : _zz_CommitPlugin_logic_reschedule_reason_2) | (_zz_CommitPlugin_logic_reschedule_reason_3 ? _zz_CommitPlugin_logic_reschedule_reason_4 : _zz_CommitPlugin_logic_reschedule_reason_5)) | ((_zz_CommitPlugin_logic_reschedule_reason_6 ? _zz_CommitPlugin_logic_reschedule_reason_7 : _zz_CommitPlugin_logic_reschedule_reason_8) | (_zz_CommitPlugin_logic_reschedule_reason_9 ? _zz_CommitPlugin_logic_reschedule_reason_10 : _zz_CommitPlugin_logic_reschedule_reason_11))) | ((CommitPlugin_logic_reschedule_portsLogic_hits[4] ? EU0_CsrAccessPlugin_setup_trap_payload_reason : 8'h00) | (CommitPlugin_logic_reschedule_portsLogic_hits[5] ? ALU1_BranchPlugin_setup_reschedule_payload_reason : 8'h00)));
      CommitPlugin_logic_reschedule_tval <= ((((CommitPlugin_logic_reschedule_portsLogic_hits[0] ? Lsu2Plugin_setup_sharedTrap_payload_tval : 32'h00000000) | (CommitPlugin_logic_reschedule_portsLogic_hits[1] ? Lsu2Plugin_setup_specialTrap_payload_tval : 32'h00000000)) | ((CommitPlugin_logic_reschedule_portsLogic_hits[2] ? ALU0_BranchPlugin_setup_reschedule_payload_tval : 32'h00000000) | (CommitPlugin_logic_reschedule_portsLogic_hits[3] ? EnvCallPlugin_setup_reschedule_payload_tval : 32'h00000000))) | ((CommitPlugin_logic_reschedule_portsLogic_hits[4] ? EU0_CsrAccessPlugin_setup_trap_payload_tval : 32'h00000000) | (CommitPlugin_logic_reschedule_portsLogic_hits[5] ? ALU1_BranchPlugin_setup_reschedule_payload_tval : 32'h00000000)));
      CommitPlugin_logic_reschedule_skipCommit <= _zz_CommitPlugin_logic_reschedule_skipCommit[0];
    end
    PrivilegedPlugin_logic_supervisor_sip_seipInput <= PrivilegedPlugin_io_int_supervisor_external;
    if(PrivilegedPlugin_logic_rescheduleUnbuffered_ready) begin
      PrivilegedPlugin_logic_rescheduleUnbuffered_rData_cause <= PrivilegedPlugin_logic_rescheduleUnbuffered_payload_cause;
      PrivilegedPlugin_logic_rescheduleUnbuffered_rData_epc <= PrivilegedPlugin_logic_rescheduleUnbuffered_payload_epc;
      PrivilegedPlugin_logic_rescheduleUnbuffered_rData_tval <= PrivilegedPlugin_logic_rescheduleUnbuffered_payload_tval;
      PrivilegedPlugin_logic_rescheduleUnbuffered_rData_fromCommit <= PrivilegedPlugin_logic_rescheduleUnbuffered_payload_fromCommit;
    end
    case(EnvCallPlugin_logic_flushes_stateReg)
      EnvCallPlugin_logic_flushes_enumDef_IDLE : begin
        if(EU0_ExecutionUnitBase_pipeline_execute_2_valid) begin
          EnvCallPlugin_logic_flushes_vmaInv <= EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA;
          EnvCallPlugin_logic_flushes_fetchInv <= EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I;
          EnvCallPlugin_logic_flushes_flushData <= EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA;
        end
      end
      EnvCallPlugin_logic_flushes_enumDef_RESCHEDULE : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_VMA_FETCH_WAIT : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_LSU_FLUSH : begin
      end
      EnvCallPlugin_logic_flushes_enumDef_WAIT_LSU : begin
      end
      default : begin
      end
    endcase
    if(Lsu2Plugin_logic_lq_regs_0_allocation) begin
      Lsu2Plugin_logic_lq_regs_0_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_0_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_1_allocation) begin
      Lsu2Plugin_logic_lq_regs_1_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_1_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_2_allocation) begin
      Lsu2Plugin_logic_lq_regs_2_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_2_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_3_allocation) begin
      Lsu2Plugin_logic_lq_regs_3_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_3_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_4_allocation) begin
      Lsu2Plugin_logic_lq_regs_4_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_4_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_5_allocation) begin
      Lsu2Plugin_logic_lq_regs_5_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_5_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_6_allocation) begin
      Lsu2Plugin_logic_lq_regs_6_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_6_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_7_allocation) begin
      Lsu2Plugin_logic_lq_regs_7_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_7_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_8_allocation) begin
      Lsu2Plugin_logic_lq_regs_8_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_8_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_9_allocation) begin
      Lsu2Plugin_logic_lq_regs_9_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_9_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_10_allocation) begin
      Lsu2Plugin_logic_lq_regs_10_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_10_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_11_allocation) begin
      Lsu2Plugin_logic_lq_regs_11_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_11_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_12_allocation) begin
      Lsu2Plugin_logic_lq_regs_12_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_12_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_13_allocation) begin
      Lsu2Plugin_logic_lq_regs_13_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_13_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_14_allocation) begin
      Lsu2Plugin_logic_lq_regs_14_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_14_niceHazard <= 1'b0;
    end
    if(Lsu2Plugin_logic_lq_regs_15_allocation) begin
      Lsu2Plugin_logic_lq_regs_15_sqChecked <= 1'b0;
      Lsu2Plugin_logic_lq_regs_15_niceHazard <= 1'b0;
    end
    Lsu2Plugin_logic_lq_ptr_priorityLast <= Lsu2Plugin_logic_lq_ptr_priority;
    Lsu2Plugin_logic_lq_tracker_freeReduced <= _zz_Lsu2Plugin_logic_lq_tracker_freeReduced;
    if(Lsu2Plugin_logic_sq_regs_0_allocation) begin
      Lsu2Plugin_logic_sq_regs_0_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_1_allocation) begin
      Lsu2Plugin_logic_sq_regs_1_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_2_allocation) begin
      Lsu2Plugin_logic_sq_regs_2_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_3_allocation) begin
      Lsu2Plugin_logic_sq_regs_3_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_4_allocation) begin
      Lsu2Plugin_logic_sq_regs_4_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_5_allocation) begin
      Lsu2Plugin_logic_sq_regs_5_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_6_allocation) begin
      Lsu2Plugin_logic_sq_regs_6_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_7_allocation) begin
      Lsu2Plugin_logic_sq_regs_7_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_8_allocation) begin
      Lsu2Plugin_logic_sq_regs_8_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_9_allocation) begin
      Lsu2Plugin_logic_sq_regs_9_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_10_allocation) begin
      Lsu2Plugin_logic_sq_regs_10_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_11_allocation) begin
      Lsu2Plugin_logic_sq_regs_11_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_12_allocation) begin
      Lsu2Plugin_logic_sq_regs_12_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_13_allocation) begin
      Lsu2Plugin_logic_sq_regs_13_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_14_allocation) begin
      Lsu2Plugin_logic_sq_regs_14_dataValid <= 1'b0;
    end
    if(Lsu2Plugin_logic_sq_regs_15_allocation) begin
      Lsu2Plugin_logic_sq_regs_15_dataValid <= 1'b0;
    end
    Lsu2Plugin_logic_sq_ptr_priorityLast <= Lsu2Plugin_logic_sq_ptr_priority;
    Lsu2Plugin_logic_sq_ptr_onFreeLast_payload <= Lsu2Plugin_logic_sq_ptr_onFree_payload;
    Lsu2Plugin_logic_sq_tracker_freeReduced <= _zz_Lsu2Plugin_logic_sq_tracker_freeReduced;
    if(Lsu2Plugin_logic_aguPush_0_pushLq) begin
      case(switch_Utils_l1437)
        4'b0000 : begin
          Lsu2Plugin_logic_lq_regs_0_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_0_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0001 : begin
          Lsu2Plugin_logic_lq_regs_1_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_1_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0010 : begin
          Lsu2Plugin_logic_lq_regs_2_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_2_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0011 : begin
          Lsu2Plugin_logic_lq_regs_3_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_3_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0100 : begin
          Lsu2Plugin_logic_lq_regs_4_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_4_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0101 : begin
          Lsu2Plugin_logic_lq_regs_5_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_5_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0110 : begin
          Lsu2Plugin_logic_lq_regs_6_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_6_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0111 : begin
          Lsu2Plugin_logic_lq_regs_7_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_7_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1000 : begin
          Lsu2Plugin_logic_lq_regs_8_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_8_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1001 : begin
          Lsu2Plugin_logic_lq_regs_9_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_9_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1010 : begin
          Lsu2Plugin_logic_lq_regs_10_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_10_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1011 : begin
          Lsu2Plugin_logic_lq_regs_11_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_11_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1100 : begin
          Lsu2Plugin_logic_lq_regs_12_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_12_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1101 : begin
          Lsu2Plugin_logic_lq_regs_13_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_13_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1110 : begin
          Lsu2Plugin_logic_lq_regs_14_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_14_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        default : begin
          Lsu2Plugin_logic_lq_regs_15_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_lq_regs_15_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
      endcase
    end
    if(when_Lsu2Plugin_l733) begin
      Lsu2Plugin_logic_sq_mem_swap <= AguPlugin_setup_port_payload_swap;
      Lsu2Plugin_logic_sq_mem_op <= AguPlugin_setup_port_payload_op;
      Lsu2Plugin_logic_sq_mem_physRd <= AguPlugin_setup_port_payload_physicalRd;
      Lsu2Plugin_logic_sq_mem_writeRd <= AguPlugin_setup_port_payload_writeRd;
    end
    if(Lsu2Plugin_logic_aguPush_0_pushSq) begin
      case(switch_Utils_l1437_1)
        4'b0000 : begin
          Lsu2Plugin_logic_sq_regs_0_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_0_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_0_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0001 : begin
          Lsu2Plugin_logic_sq_regs_1_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_1_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_1_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0010 : begin
          Lsu2Plugin_logic_sq_regs_2_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_2_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_2_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0011 : begin
          Lsu2Plugin_logic_sq_regs_3_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_3_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_3_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0100 : begin
          Lsu2Plugin_logic_sq_regs_4_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_4_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_4_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0101 : begin
          Lsu2Plugin_logic_sq_regs_5_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_5_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_5_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0110 : begin
          Lsu2Plugin_logic_sq_regs_6_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_6_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_6_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b0111 : begin
          Lsu2Plugin_logic_sq_regs_7_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_7_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_7_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1000 : begin
          Lsu2Plugin_logic_sq_regs_8_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_8_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_8_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1001 : begin
          Lsu2Plugin_logic_sq_regs_9_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_9_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_9_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1010 : begin
          Lsu2Plugin_logic_sq_regs_10_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_10_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_10_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1011 : begin
          Lsu2Plugin_logic_sq_regs_11_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_11_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_11_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1100 : begin
          Lsu2Plugin_logic_sq_regs_12_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_12_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_12_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1101 : begin
          Lsu2Plugin_logic_sq_regs_13_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_13_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_13_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        4'b1110 : begin
          Lsu2Plugin_logic_sq_regs_14_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_14_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_14_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
        default : begin
          Lsu2Plugin_logic_sq_regs_15_dataValid <= 1'b1;
          Lsu2Plugin_logic_sq_regs_15_address_pageOffset <= AguPlugin_setup_port_payload_address[11 : 2];
          Lsu2Plugin_logic_sq_regs_15_address_mask <= Lsu2Plugin_logic_aguPush_0_dataMask;
        end
      endcase
    end
    if(when_Lsu2Plugin_l1046) begin
      case(Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID)
        4'b0000 : begin
          Lsu2Plugin_logic_lq_regs_0_sqChecked <= 1'b1;
        end
        4'b0001 : begin
          Lsu2Plugin_logic_lq_regs_1_sqChecked <= 1'b1;
        end
        4'b0010 : begin
          Lsu2Plugin_logic_lq_regs_2_sqChecked <= 1'b1;
        end
        4'b0011 : begin
          Lsu2Plugin_logic_lq_regs_3_sqChecked <= 1'b1;
        end
        4'b0100 : begin
          Lsu2Plugin_logic_lq_regs_4_sqChecked <= 1'b1;
        end
        4'b0101 : begin
          Lsu2Plugin_logic_lq_regs_5_sqChecked <= 1'b1;
        end
        4'b0110 : begin
          Lsu2Plugin_logic_lq_regs_6_sqChecked <= 1'b1;
        end
        4'b0111 : begin
          Lsu2Plugin_logic_lq_regs_7_sqChecked <= 1'b1;
        end
        4'b1000 : begin
          Lsu2Plugin_logic_lq_regs_8_sqChecked <= 1'b1;
        end
        4'b1001 : begin
          Lsu2Plugin_logic_lq_regs_9_sqChecked <= 1'b1;
        end
        4'b1010 : begin
          Lsu2Plugin_logic_lq_regs_10_sqChecked <= 1'b1;
        end
        4'b1011 : begin
          Lsu2Plugin_logic_lq_regs_11_sqChecked <= 1'b1;
        end
        4'b1100 : begin
          Lsu2Plugin_logic_lq_regs_12_sqChecked <= 1'b1;
        end
        4'b1101 : begin
          Lsu2Plugin_logic_lq_regs_13_sqChecked <= 1'b1;
        end
        4'b1110 : begin
          Lsu2Plugin_logic_lq_regs_14_sqChecked <= 1'b1;
        end
        default : begin
          Lsu2Plugin_logic_lq_regs_15_sqChecked <= 1'b1;
        end
      endcase
    end
    if(when_Lsu2Plugin_l1104) begin
      Lsu2Plugin_logic_lq_regs_0_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_1) begin
      Lsu2Plugin_logic_lq_regs_1_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_2) begin
      Lsu2Plugin_logic_lq_regs_2_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_3) begin
      Lsu2Plugin_logic_lq_regs_3_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_4) begin
      Lsu2Plugin_logic_lq_regs_4_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_5) begin
      Lsu2Plugin_logic_lq_regs_5_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_6) begin
      Lsu2Plugin_logic_lq_regs_6_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_7) begin
      Lsu2Plugin_logic_lq_regs_7_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_8) begin
      Lsu2Plugin_logic_lq_regs_8_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_9) begin
      Lsu2Plugin_logic_lq_regs_9_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_10) begin
      Lsu2Plugin_logic_lq_regs_10_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_11) begin
      Lsu2Plugin_logic_lq_regs_11_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_12) begin
      Lsu2Plugin_logic_lq_regs_12_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_13) begin
      Lsu2Plugin_logic_lq_regs_13_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_14) begin
      Lsu2Plugin_logic_lq_regs_14_niceHazard <= 1'b1;
    end
    if(when_Lsu2Plugin_l1104_15) begin
      Lsu2Plugin_logic_lq_regs_15_niceHazard <= 1'b1;
    end
    if(Lsu2Plugin_logic_sharedPip_stages_3_isFireing) begin
      case(Lsu2Plugin_logic_sharedPip_stages_3_CTRL)
        Lsu2Plugin_CTRL_ENUM_TRAP_ALIGN : begin
        end
        Lsu2Plugin_CTRL_ENUM_MMU_REDO : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_MMU : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_HAZARD : begin
          if(_zz_103) begin
            Lsu2Plugin_logic_lq_regs_0_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_104) begin
            Lsu2Plugin_logic_lq_regs_1_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_105) begin
            Lsu2Plugin_logic_lq_regs_2_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_106) begin
            Lsu2Plugin_logic_lq_regs_3_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_107) begin
            Lsu2Plugin_logic_lq_regs_4_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_108) begin
            Lsu2Plugin_logic_lq_regs_5_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_109) begin
            Lsu2Plugin_logic_lq_regs_6_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_110) begin
            Lsu2Plugin_logic_lq_regs_7_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_111) begin
            Lsu2Plugin_logic_lq_regs_8_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_112) begin
            Lsu2Plugin_logic_lq_regs_9_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_113) begin
            Lsu2Plugin_logic_lq_regs_10_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_114) begin
            Lsu2Plugin_logic_lq_regs_11_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_115) begin
            Lsu2Plugin_logic_lq_regs_12_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_116) begin
            Lsu2Plugin_logic_lq_regs_13_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_117) begin
            Lsu2Plugin_logic_lq_regs_14_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
          if(_zz_118) begin
            Lsu2Plugin_logic_lq_regs_15_waitOn_sqId <= _zz_Lsu2Plugin_logic_lq_regs_0_waitOn_sqId;
          end
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_MISS : begin
        end
        Lsu2Plugin_CTRL_ENUM_LOAD_FAILED : begin
        end
        Lsu2Plugin_CTRL_ENUM_TRAP_ACCESS : begin
        end
        default : begin
          if(Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD) begin
            if(when_Lsu2Plugin_l1333) begin
              if(Lsu2Plugin_logic_sharedPip_stages_3_LR) begin
                Lsu2Plugin_logic_lq_reservation_address <= Lsu2Plugin_logic_sharedPip_stages_3_MMU_TRANSLATED;
              end
            end
          end
        end
      endcase
    end
    if(Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_ready) begin
      toplevel_Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_rData <= Lsu2Plugin_logic_prefetch_predictor_io_prediction_cmd_payload;
    end
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_fault <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_fault;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_redo <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_redo;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlot <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlot;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_refillSlotAny <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_refillSlotAny;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_generationKo <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_generationKo;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_flush <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_flush;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_prefetch <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_prefetch;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_address <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_address;
    Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_regNext_payload_io <= Lsu2Plugin_logic_writeback_rsp_delayed_0_combStage_payload_io;
    if(Lsu2Plugin_setup_flushPort_cmd_valid) begin
      Lsu2Plugin_logic_flush_cmdPtr <= 7'h00;
      Lsu2Plugin_logic_flush_rspPtr <= 7'h00;
      Lsu2Plugin_logic_flush_withFree <= Lsu2Plugin_setup_flushPort_cmd_payload_withFree;
    end
    if(when_Lsu2Plugin_l1553) begin
      if(Lsu2Plugin_setup_cacheStore_cmd_fire) begin
        Lsu2Plugin_logic_flush_cmdPtr <= (Lsu2Plugin_logic_flush_cmdPtr + 7'h01);
      end
      if(when_Lsu2Plugin_l1561) begin
        if(Lsu2Plugin_setup_cacheStore_rsp_payload_redo) begin
          Lsu2Plugin_logic_flush_cmdPtr <= Lsu2Plugin_logic_flush_rspPtr;
        end else begin
          Lsu2Plugin_logic_flush_rspPtr <= (Lsu2Plugin_logic_flush_rspPtr + 7'h01);
        end
      end
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_isStore <= Lsu2Plugin_logic_special_storeHit;
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_isLoad <= (! Lsu2Plugin_logic_special_storeHit);
    end
    Lsu2Plugin_logic_special_robId <= CommitPlugin_logic_commit_head;
    Lsu2Plugin_logic_special_loadPhysRd <= _zz_Lsu2Plugin_logic_lq_mem_physRd_port2;
    Lsu2Plugin_logic_special_loadAddress <= _zz_Lsu2Plugin_logic_lq_mem_addressPost_port2;
    Lsu2Plugin_logic_special_loadAddressVirt <= _zz_Lsu2Plugin_logic_lq_mem_addressPre_port2;
    Lsu2Plugin_logic_special_loadSize <= _zz_Lsu2Plugin_logic_lq_mem_size_port2;
    Lsu2Plugin_logic_special_loadUnsigned <= _zz_Lsu2Plugin_logic_lq_mem_unsigned_port2[0];
    Lsu2Plugin_logic_special_loadWriteRd <= (Lsu2Plugin_logic_special_isLoad && _zz_Lsu2Plugin_logic_lq_mem_writeRd_port2[0]);
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeAddress <= Lsu2Plugin_setup_cacheStore_cmd_payload_address;
    end
    Lsu2Plugin_logic_special_storeAddressVirt <= _zz_Lsu2Plugin_logic_sq_mem_addressPre_port2;
    Lsu2Plugin_logic_special_storeSize <= _zz_Lsu2Plugin_logic_sq_mem_size_port4;
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeData <= Lsu2Plugin_setup_cacheStore_cmd_payload_data;
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeMask <= Lsu2Plugin_setup_cacheStore_cmd_payload_mask;
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeAmo <= _zz_Lsu2Plugin_logic_sq_mem_amo_port2[0];
    end
    if(Lsu2Plugin_logic_special_hit) begin
      Lsu2Plugin_logic_special_storeSc <= _zz_Lsu2Plugin_logic_sq_mem_sc_port2[0];
    end
    if(PrivilegedPlugin_logic_decoderInterrupt_buffer_sample) begin
      PrivilegedPlugin_logic_decoderInterrupt_buffer_code <= PrivilegedPlugin_logic_interrupt_code;
    end
    if(PrivilegedPlugin_logic_decoderInterrupt_buffer_sample) begin
      PrivilegedPlugin_logic_decoderInterrupt_buffer_targetPrivilege <= PrivilegedPlugin_logic_interrupt_targetPrivilege;
    end
    MmuPlugin_logic_refill_portsOh_regNext <= MmuPlugin_logic_refill_portsOh;
    _zz_MmuPlugin_logic_refill_portsAddress <= Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION;
    _zz_MmuPlugin_logic_refill_portsAddress_1 <= FetchPlugin_stages_1_Fetch_FETCH_PC;
    MmuPlugin_logic_refill_load_rsp_payload_data <= MmuPlugin_setup_cacheLoad_rsp_payload_data;
    MmuPlugin_logic_refill_load_rsp_payload_fault <= MmuPlugin_setup_cacheLoad_rsp_payload_fault;
    MmuPlugin_logic_refill_load_rsp_payload_redo <= MmuPlugin_setup_cacheLoad_rsp_payload_redo;
    MmuPlugin_logic_refill_load_rsp_payload_refillSlot <= MmuPlugin_setup_cacheLoad_rsp_payload_refillSlot;
    MmuPlugin_logic_refill_load_rsp_payload_refillSlotAny <= MmuPlugin_setup_cacheLoad_rsp_payload_refillSlotAny;
    Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION <= Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION;
    Lsu2Plugin_logic_sharedPip_stages_1_ROB_ID <= Lsu2Plugin_logic_sharedPip_stages_0_ROB_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_PHYS_RD <= Lsu2Plugin_logic_sharedPip_stages_0_PHYS_RD;
    Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_PRE_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_POST_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_0_ADDRESS_POST_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_1_SIZE <= Lsu2Plugin_logic_sharedPip_stages_0_SIZE;
    Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_0_NEED_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_1_TRANSLATED_AS_IO <= Lsu2Plugin_logic_sharedPip_stages_0_TRANSLATED_AS_IO;
    Lsu2Plugin_logic_sharedPip_stages_1_WRITE_RD <= Lsu2Plugin_logic_sharedPip_stages_0_WRITE_RD;
    Lsu2Plugin_logic_sharedPip_stages_1_UNSIGNED <= Lsu2Plugin_logic_sharedPip_stages_0_UNSIGNED;
    Lsu2Plugin_logic_sharedPip_stages_1_LR <= Lsu2Plugin_logic_sharedPip_stages_0_LR;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_VALID <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_VALID;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_DELTA <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_DELTA;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SCORE <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SCORE;
    Lsu2Plugin_logic_sharedPip_stages_1_AMO <= Lsu2Plugin_logic_sharedPip_stages_0_AMO;
    Lsu2Plugin_logic_sharedPip_stages_1_SC <= Lsu2Plugin_logic_sharedPip_stages_0_SC;
    Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD <= Lsu2Plugin_logic_sharedPip_stages_0_IS_LOAD;
    Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID <= Lsu2Plugin_logic_sharedPip_stages_0_LQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID <= Lsu2Plugin_logic_sharedPip_stages_0_SQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH;
    Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION_COUNTER <= Lsu2Plugin_logic_sharedPip_stages_0_HIT_SPECULATION_COUNTER;
    Lsu2Plugin_logic_sharedPip_stages_1_SP_FP_ADDRESS <= Lsu2Plugin_logic_sharedPip_stages_0_SP_FP_ADDRESS;
    Lsu2Plugin_logic_sharedPip_stages_1_DATA_MASK <= Lsu2Plugin_logic_sharedPip_stages_0_DATA_MASK;
    Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_START_ID <= Lsu2Plugin_logic_sharedPip_stages_0_LQCHECK_START_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_SQCHECK_END_ID <= Lsu2Plugin_logic_sharedPip_stages_0_SQCHECK_END_ID;
    Lsu2Plugin_logic_sharedPip_stages_1_feed_SQ_PTR_FREE <= Lsu2Plugin_logic_sharedPip_stages_0_feed_SQ_PTR_FREE;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SQID <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_SQID;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_HAZARD_PRED_HIT_FEEDED;
    Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH_PC <= Lsu2Plugin_logic_sharedPip_stages_0_LOAD_FRESH_PC;
    Lsu2Plugin_logic_sharedPip_stages_1_MmuPlugin_logic_ALLOW_REFILL <= Lsu2Plugin_logic_sharedPip_stages_0_MmuPlugin_logic_ALLOW_REFILL_overloaded;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_0_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_0_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_1_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_1_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_2_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_2_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_ENTRIES_3_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_ENTRIES_3_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L0_HITS_PRE_VALID <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L0_HITS_PRE_VALID;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_0_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_0_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_valid <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_valid;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_pageFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_pageFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_accessFault <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_accessFault;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_virtualAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_virtualAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_physicalAddress <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_physicalAddress;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowRead <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowRead;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowWrite <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowWrite;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowExecute <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowExecute;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_ENTRIES_1_allowUser <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_ENTRIES_1_allowUser;
    Lsu2Plugin_logic_sharedPip_stages_1_MMU_L1_HITS_PRE_VALID <= Lsu2Plugin_logic_sharedPip_stages_0_MMU_L1_HITS_PRE_VALID;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SQID <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SQID;
    Lsu2Plugin_logic_sharedPip_stages_2_NEED_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_1_NEED_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_TRANSLATED <= Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_TRANSLATED;
    Lsu2Plugin_logic_sharedPip_stages_2_IS_IO <= Lsu2Plugin_logic_sharedPip_stages_1_IS_IO;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_TRANSLATED <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_TRANSLATED;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_PAGE_FAULT <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_PAGE_FAULT;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_ACCESS_FAULT <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_ACCESS_FAULT;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_READ <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_READ;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_REDO <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_REDO;
    Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_1_ADDRESS_PRE_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_HIT <= Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_HIT;
    Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID <= Lsu2Plugin_logic_sharedPip_stages_1_OLDER_STORE_ID;
    Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD <= Lsu2Plugin_logic_sharedPip_stages_1_IS_LOAD;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_HIT;
    Lsu2Plugin_logic_sharedPip_stages_2_LQ_ID <= Lsu2Plugin_logic_sharedPip_stages_1_LQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_2_SQ_ID <= Lsu2Plugin_logic_sharedPip_stages_1_SQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_HITS <= Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_HITS;
    Lsu2Plugin_logic_sharedPip_stages_2_LQCHECK_NO_YOUNGER <= Lsu2Plugin_logic_sharedPip_stages_1_LQCHECK_NO_YOUNGER;
    Lsu2Plugin_logic_sharedPip_stages_2_MMU_ALLOW_WRITE <= Lsu2Plugin_logic_sharedPip_stages_1_MMU_ALLOW_WRITE;
    Lsu2Plugin_logic_sharedPip_stages_2_SIZE <= Lsu2Plugin_logic_sharedPip_stages_1_SIZE;
    Lsu2Plugin_logic_sharedPip_stages_2_UNSIGNED <= Lsu2Plugin_logic_sharedPip_stages_1_UNSIGNED;
    Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID <= Lsu2Plugin_logic_sharedPip_stages_1_ROB_ID;
    Lsu2Plugin_logic_sharedPip_stages_2_WRITE_RD <= Lsu2Plugin_logic_sharedPip_stages_1_WRITE_RD;
    Lsu2Plugin_logic_sharedPip_stages_2_PHYS_RD <= Lsu2Plugin_logic_sharedPip_stages_1_PHYS_RD;
    Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION <= Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION;
    Lsu2Plugin_logic_sharedPip_stages_2_LR <= Lsu2Plugin_logic_sharedPip_stages_1_LR;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SCORE <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_SCORE;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_VALID <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_VALID;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_DELTA <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_HAZARD_PRED_DELTA;
    Lsu2Plugin_logic_sharedPip_stages_2_SC <= Lsu2Plugin_logic_sharedPip_stages_1_SC;
    Lsu2Plugin_logic_sharedPip_stages_2_AMO <= Lsu2Plugin_logic_sharedPip_stages_1_AMO;
    Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION_COUNTER <= Lsu2Plugin_logic_sharedPip_stages_1_HIT_SPECULATION_COUNTER;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH;
    Lsu2Plugin_logic_sharedPip_stages_2_SP_FP_ADDRESS <= Lsu2Plugin_logic_sharedPip_stages_1_SP_FP_ADDRESS;
    Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH_PC <= Lsu2Plugin_logic_sharedPip_stages_1_LOAD_FRESH_PC;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT_FEEDED <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT_FEEDED_overloaded;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SQID <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SQID;
    Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_COMPLETED <= Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_COMPLETED_overloaded;
    Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_ID <= Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_OLDER_STORE_WAIT_FEED <= Lsu2Plugin_logic_sharedPip_stages_2_OLDER_STORE_WAIT_FEED;
    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ROB <= Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ROB;
    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_RESCHEDULE <= Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_RESCHEDULE;
    Lsu2Plugin_logic_sharedPip_stages_3_YOUNGER_LOAD_ID <= Lsu2Plugin_logic_sharedPip_stages_2_YOUNGER_LOAD_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_valid <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_valid;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_data <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_data;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_fault <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_fault;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_redo <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_redo;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlot <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlot;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_CACHE_RSP_payload_refillSlotAny <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_CACHE_RSP_overloaded_payload_refillSlotAny;
    Lsu2Plugin_logic_sharedPip_stages_3_ADDRESS_PRE_TRANSLATION <= Lsu2Plugin_logic_sharedPip_stages_2_ADDRESS_PRE_TRANSLATION;
    Lsu2Plugin_logic_sharedPip_stages_3_IS_IO <= Lsu2Plugin_logic_sharedPip_stages_2_IS_IO;
    Lsu2Plugin_logic_sharedPip_stages_3_IS_LOAD <= Lsu2Plugin_logic_sharedPip_stages_2_IS_LOAD;
    Lsu2Plugin_logic_sharedPip_stages_3_ROB_ID <= Lsu2Plugin_logic_sharedPip_stages_2_ROB_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_LQ_ID <= Lsu2Plugin_logic_sharedPip_stages_2_LQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_WRITE_RD <= Lsu2Plugin_logic_sharedPip_stages_2_WRITE_RD;
    Lsu2Plugin_logic_sharedPip_stages_3_PHYS_RD <= Lsu2Plugin_logic_sharedPip_stages_2_PHYS_RD;
    Lsu2Plugin_logic_sharedPip_stages_3_CTRL <= Lsu2Plugin_logic_sharedPip_stages_2_CTRL;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_HIT <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_HIT;
    Lsu2Plugin_logic_sharedPip_stages_3_TRAP_SPECULATION <= Lsu2Plugin_logic_sharedPip_stages_2_TRAP_SPECULATION;
    Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION <= Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION;
    Lsu2Plugin_logic_sharedPip_stages_3_SQ_ID <= Lsu2Plugin_logic_sharedPip_stages_2_SQ_ID;
    Lsu2Plugin_logic_sharedPip_stages_3_LR <= Lsu2Plugin_logic_sharedPip_stages_2_LR;
    Lsu2Plugin_logic_sharedPip_stages_3_MMU_TRANSLATED <= Lsu2Plugin_logic_sharedPip_stages_2_MMU_TRANSLATED;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_SCORE <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_SCORE;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_VALID <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_VALID;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_HAZARD_PRED_DELTA <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_HAZARD_PRED_DELTA;
    Lsu2Plugin_logic_sharedPip_stages_3_SC <= Lsu2Plugin_logic_sharedPip_stages_2_SC;
    Lsu2Plugin_logic_sharedPip_stages_3_AMO <= Lsu2Plugin_logic_sharedPip_stages_2_AMO;
    Lsu2Plugin_logic_sharedPip_stages_3_HIT_SPECULATION_COUNTER <= Lsu2Plugin_logic_sharedPip_stages_2_HIT_SPECULATION_COUNTER;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH;
    Lsu2Plugin_logic_sharedPip_stages_3_SP_FP_ADDRESS <= Lsu2Plugin_logic_sharedPip_stages_2_SP_FP_ADDRESS;
    Lsu2Plugin_logic_sharedPip_stages_3_LOAD_FRESH_PC <= Lsu2Plugin_logic_sharedPip_stages_2_LOAD_FRESH_PC;
    if(Lsu2Plugin_logic_lqSqArbitration_s0_ready_output) begin
      Lsu2Plugin_logic_lqSqArbitration_s1_LQ_HIT <= Lsu2Plugin_logic_lqSqArbitration_s0_LQ_HIT;
      Lsu2Plugin_logic_lqSqArbitration_s1_SQ_HIT <= Lsu2Plugin_logic_lqSqArbitration_s0_SQ_HIT;
      Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ID <= Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ID;
      Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ID <= Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ID;
      Lsu2Plugin_logic_lqSqArbitration_s1_LQ_ROB_FULL <= Lsu2Plugin_logic_lqSqArbitration_s0_LQ_ROB_FULL;
      Lsu2Plugin_logic_lqSqArbitration_s1_SQ_ROB_FULL <= Lsu2Plugin_logic_lqSqArbitration_s0_SQ_ROB_FULL;
    end
    (* parallel_case *)
    case(1) // synthesis parallel_case
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_IDLE) == Lsu2Plugin_logic_special_atomic_enumDef_IDLE) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_CMD) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) == Lsu2Plugin_logic_special_atomic_enumDef_LOAD_RSP) : begin
        Lsu2Plugin_logic_special_atomic_readed <= Lsu2Plugin_logic_sharedPip_cacheRsp_rspFormated[31 : 0];
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) == Lsu2Plugin_logic_special_atomic_enumDef_LOCK_DELAY) : begin
        if(when_Lsu2Plugin_l1715) begin
          Lsu2Plugin_logic_special_atomic_gotReservation <= (Lsu2Plugin_logic_lq_reservation_valid && (Lsu2Plugin_logic_lq_reservation_address == Lsu2Plugin_logic_special_storeAddress));
        end
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_ALU) == Lsu2Plugin_logic_special_atomic_enumDef_ALU) : begin
        Lsu2Plugin_logic_special_atomic_result <= Lsu2Plugin_logic_special_atomic_alu_result;
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) == Lsu2Plugin_logic_special_atomic_enumDef_COMPLETION) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_SYNC) == Lsu2Plugin_logic_special_atomic_enumDef_SYNC) : begin
      end
      (((Lsu2Plugin_logic_special_atomic_stateReg) & Lsu2Plugin_logic_special_atomic_enumDef_TRAP) == Lsu2Plugin_logic_special_atomic_enumDef_TRAP) : begin
      end
      default : begin
      end
    endcase
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_enumDef_IDLE : begin
        MmuPlugin_logic_refill_portOhReg <= MmuPlugin_logic_refill_portsOh;
      end
      MmuPlugin_logic_refill_enumDef_INIT : begin
        MmuPlugin_logic_refill_virtual <= MmuPlugin_logic_refill_portsAddress;
        MmuPlugin_logic_refill_load_address <= {{MmuPlugin_logic_satp_ppn,MmuPlugin_logic_refill_portsAddress[31 : 22]},2'b00};
      end
      MmuPlugin_logic_refill_enumDef_CMD_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_CMD_1 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_0 : begin
      end
      MmuPlugin_logic_refill_enumDef_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(!when_MmuPlugin_l469) begin
              MmuPlugin_logic_refill_load_address <= MmuPlugin_logic_refill_load_nextLevelBase;
              MmuPlugin_logic_refill_load_address[11 : 2] <= MmuPlugin_logic_refill_virtual[21 : 12];
            end
          end
        end
      end
      default : begin
      end
    endcase
    case(EU0_CsrAccessPlugin_logic_fsm_stateReg)
      EU0_CsrAccessPlugin_logic_fsm_enumDef_IDLE : begin
        EU0_CsrAccessPlugin_logic_fsm_regs_microOp <= EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
        EU0_CsrAccessPlugin_logic_fsm_regs_doImm <= EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_IMM;
        EU0_CsrAccessPlugin_logic_fsm_regs_doMask <= EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_MASK;
        EU0_CsrAccessPlugin_logic_fsm_regs_doClear <= EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_CSR_CLEAR;
        EU0_CsrAccessPlugin_logic_fsm_regs_rs1 <= EU0_ExecutionUnitBase_pipeline_execute_0_integer_RS1;
        EU0_CsrAccessPlugin_logic_fsm_regs_implemented <= EU0_CsrAccessPlugin_logic_fsm_startLogic_implemented;
        EU0_CsrAccessPlugin_logic_fsm_regs_trap <= EU0_CsrAccessPlugin_logic_fsm_startLogic_trap;
        EU0_CsrAccessPlugin_logic_fsm_regs_flushPipeline <= EU0_CsrAccessPlugin_setup_onDecodeFlushPipeline;
        EU0_CsrAccessPlugin_logic_fsm_regs_write <= EU0_CsrAccessPlugin_logic_fsm_startLogic_write;
        EU0_CsrAccessPlugin_logic_fsm_regs_read <= EU0_CsrAccessPlugin_logic_fsm_startLogic_read;
        REG_CSR_773 <= COMB_CSR_773;
        REG_CSR_835 <= COMB_CSR_835;
        REG_CSR_833 <= COMB_CSR_833;
        REG_CSR_832 <= COMB_CSR_832;
        REG_CSR_3857 <= COMB_CSR_3857;
        REG_CSR_3858 <= COMB_CSR_3858;
        REG_CSR_3859 <= COMB_CSR_3859;
        REG_CSR_3860 <= COMB_CSR_3860;
        REG_CSR_769 <= COMB_CSR_769;
        REG_CSR_834 <= COMB_CSR_834;
        REG_CSR_768 <= COMB_CSR_768;
        REG_CSR_836 <= COMB_CSR_836;
        REG_CSR_772 <= COMB_CSR_772;
        REG_CSR_770 <= COMB_CSR_770;
        REG_CSR_771 <= COMB_CSR_771;
        REG_CSR_261 <= COMB_CSR_261;
        REG_CSR_323 <= COMB_CSR_323;
        REG_CSR_321 <= COMB_CSR_321;
        REG_CSR_320 <= COMB_CSR_320;
        REG_CSR_322 <= COMB_CSR_322;
        REG_CSR_256 <= COMB_CSR_256;
        REG_CSR_260 <= COMB_CSR_260;
        REG_CSR_324 <= COMB_CSR_324;
        REG_CSR_262 <= COMB_CSR_262;
        REG_CSR_774 <= COMB_CSR_774;
        REG_CSR_ <= COMB_CSR_;
        REG_CSR_803 <= COMB_CSR_803;
        REG_CSR_804 <= COMB_CSR_804;
        REG_CSR_805 <= COMB_CSR_805;
        REG_CSR_806 <= COMB_CSR_806;
        REG_CSR_384 <= COMB_CSR_384;
        REG_CSR_PerformanceCounterPlugin_logic_csrFilter <= COMB_CSR_PerformanceCounterPlugin_logic_csrFilter;
        EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b0;
        case(switch_CsrAccessPlugin_l204)
          12'h305 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 5'h17;
          end
          12'h343 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 5'h16;
          end
          12'h341 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 5'h15;
          end
          12'h340 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 5'h14;
          end
          12'h105 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 5'h13;
          end
          12'h143 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 5'h12;
          end
          12'h141 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 5'h11;
          end
          12'h140 : begin
            EU0_CsrAccessPlugin_logic_fsm_regs_ramSel <= 1'b1;
            EU0_CsrAccessPlugin_logic_fsm_regs_ramAddress <= 5'h10;
          end
          default : begin
          end
        endcase
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_READ : begin
        EU0_CsrAccessPlugin_logic_fsm_regs_aluInput <= EU0_CsrAccessPlugin_setup_onReadToWriteBits;
        EU0_CsrAccessPlugin_logic_fsm_regs_csrValue <= EU0_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_WRITE : begin
        if(EU0_CsrAccessPlugin_setup_onWriteFlushPipeline) begin
          EU0_CsrAccessPlugin_logic_fsm_regs_flushPipeline <= 1'b1;
        end
      end
      EU0_CsrAccessPlugin_logic_fsm_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
    if(when_DecoderPlugin_l302) begin
      DecoderPlugin_logic_exception_exceptionReg_0 <= FrontendPlugin_decoded_TRAP_0;
      DecoderPlugin_logic_exception_exceptionReg_1 <= FrontendPlugin_decoded_TRAP_1;
    end
    if(when_DecoderPlugin_l303) begin
      DecoderPlugin_logic_exception_fetchFaultReg_0 <= FrontendPlugin_decoded_Frontend_FETCH_FAULT_0;
      DecoderPlugin_logic_exception_fetchFaultReg_1 <= FrontendPlugin_decoded_Frontend_FETCH_FAULT_1;
    end
    if(when_DecoderPlugin_l304) begin
      DecoderPlugin_logic_exception_fetchFaultPageReg_0 <= FrontendPlugin_decoded_Frontend_FETCH_FAULT_PAGE_0;
      DecoderPlugin_logic_exception_fetchFaultPageReg_1 <= FrontendPlugin_decoded_Frontend_FETCH_FAULT_PAGE_1;
    end
    if(when_DecoderPlugin_l306) begin
      DecoderPlugin_logic_exception_debugEnterReg_0 <= DecoderPlugin_setup_debugEnter_0;
      DecoderPlugin_logic_exception_debugEnterReg_1 <= DecoderPlugin_setup_debugEnter_1;
    end
    if(when_DecoderPlugin_l307) begin
      DecoderPlugin_logic_exception_epcReg_0 <= FrontendPlugin_decoded_PC_0;
      DecoderPlugin_logic_exception_epcReg_1 <= FrontendPlugin_decoded_PC_1;
    end
    if(when_DecoderPlugin_l308) begin
      DecoderPlugin_logic_exception_instReg_0 <= FrontendPlugin_decoded_Frontend_INSTRUCTION_ALIGNED_0;
      DecoderPlugin_logic_exception_instReg_1 <= FrontendPlugin_decoded_Frontend_INSTRUCTION_ALIGNED_1;
    end
    ALU0_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP <= ALU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1 <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2 <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_PC <= ALU0_ExecutionUnitBase_pipeline_fetch_0_PC;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID <= ALU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD <= ALU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD <= ALU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_BRANCH_ID <= ALU0_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_SEL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E0 <= ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SEL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_LEFT <= ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SIGNED <= ALU0_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_SEL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E1 <= ALU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL <= ALU0_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
    ALU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED <= ALU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
    ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL <= ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL;
    ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND <= ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
    ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL <= ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL;
    ALU0_ExecutionUnitBase_pipeline_execute_1_PC <= ALU0_ExecutionUnitBase_pipeline_execute_0_PC;
    ALU0_ExecutionUnitBase_pipeline_execute_1_PC_TRUE <= ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TRUE;
    ALU0_ExecutionUnitBase_pipeline_execute_1_PC_TARGET <= ALU0_ExecutionUnitBase_pipeline_execute_0_PC_TARGET;
    ALU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_taken <= ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken;
    ALU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_pc <= ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc;
    ALU0_ExecutionUnitBase_pipeline_execute_1_BRANCH_ID <= ALU0_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID;
    ALU0_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BAD_EARLY_TARGET <= ALU0_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BAD_EARLY_TARGET;
    ALU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID <= ALU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
    ALU0_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E1 <= ALU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E1;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP <= ALU1_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1 <= ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2 <= ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_PC <= ALU1_ExecutionUnitBase_pipeline_fetch_0_PC;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_ROB_ID <= ALU1_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD <= ALU1_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD <= ALU1_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_BRANCH_ID <= ALU1_ExecutionUnitBase_pipeline_fetch_0_BRANCH_ID;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_SEL <= ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_SEL;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E0 <= ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E0;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_CTRL <= ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_CTRL;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_IntAluPlugin_ALU_BITWISE_CTRL <= ALU1_ExecutionUnitBase_pipeline_fetch_0_IntAluPlugin_ALU_BITWISE_CTRL;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SEL <= ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SEL;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_LEFT <= ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_LEFT;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_ShiftPlugin_SIGNED <= ALU1_ExecutionUnitBase_pipeline_fetch_0_ShiftPlugin_SIGNED;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_SEL <= ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_SEL;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E1 <= ALU1_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E1;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_BranchPlugin_BRANCH_CTRL <= ALU1_ExecutionUnitBase_pipeline_fetch_0_BranchPlugin_BRANCH_CTRL;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT <= ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO <= ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
    ALU1_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_UNSIGNED <= ALU1_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_UNSIGNED;
    ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_SEL <= ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_SEL;
    ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_COND <= ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_COND;
    ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BRANCH_CTRL <= ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BRANCH_CTRL;
    ALU1_ExecutionUnitBase_pipeline_execute_1_PC <= ALU1_ExecutionUnitBase_pipeline_execute_0_PC;
    ALU1_ExecutionUnitBase_pipeline_execute_1_PC_TRUE <= ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TRUE;
    ALU1_ExecutionUnitBase_pipeline_execute_1_PC_TARGET <= ALU1_ExecutionUnitBase_pipeline_execute_0_PC_TARGET;
    ALU1_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_taken <= ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_taken;
    ALU1_ExecutionUnitBase_pipeline_execute_1_BRANCH_EARLY_pc <= ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_EARLY_pc;
    ALU1_ExecutionUnitBase_pipeline_execute_1_BRANCH_ID <= ALU1_ExecutionUnitBase_pipeline_execute_0_BRANCH_ID;
    ALU1_ExecutionUnitBase_pipeline_execute_1_BranchPlugin_BAD_EARLY_TARGET <= ALU1_ExecutionUnitBase_pipeline_execute_0_BranchPlugin_BAD_EARLY_TARGET;
    ALU1_ExecutionUnitBase_pipeline_execute_1_ROB_ID <= ALU1_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
    ALU1_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E1 <= ALU1_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E1;
    if(EU0_ExecutionUnitBase_pipeline_fetch_0_ready_output) begin
      EU0_ExecutionUnitBase_pipeline_fetch_1_Frontend_MICRO_OP <= EU0_ExecutionUnitBase_pipeline_fetch_0_Frontend_MICRO_OP;
      EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC1 <= EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC1;
      EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS1 <= EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS1;
      EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_SRC2 <= EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_SRC2;
      EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_ID <= EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_ID;
      EU0_ExecutionUnitBase_pipeline_fetch_1_PHYS_RD <= EU0_ExecutionUnitBase_pipeline_fetch_0_PHYS_RD;
      EU0_ExecutionUnitBase_pipeline_fetch_1_WRITE_RD <= EU0_ExecutionUnitBase_pipeline_fetch_0_WRITE_RD;
      EU0_ExecutionUnitBase_pipeline_fetch_1_PC <= EU0_ExecutionUnitBase_pipeline_fetch_0_PC;
      EU0_ExecutionUnitBase_pipeline_fetch_1_LSU_ID <= EU0_ExecutionUnitBase_pipeline_fetch_0_LSU_ID;
      EU0_ExecutionUnitBase_pipeline_fetch_1_ROB_MSB <= EU0_ExecutionUnitBase_pipeline_fetch_0_ROB_MSB;
      EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_completion_SEL_E2 <= EU0_ExecutionUnitBase_pipeline_fetch_0_completion_SEL_E2;
      EU0_ExecutionUnitBase_pipeline_fetch_1_MulPlugin_HIGH <= EU0_ExecutionUnitBase_pipeline_fetch_0_MulPlugin_HIGH;
      EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS1_SIGNED <= EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS1_SIGNED;
      EU0_ExecutionUnitBase_pipeline_fetch_1_RsUnsignedPlugin_RS2_SIGNED <= EU0_ExecutionUnitBase_pipeline_fetch_0_RsUnsignedPlugin_RS2_SIGNED;
      EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_DivPlugin_REM <= EU0_ExecutionUnitBase_pipeline_fetch_0_DivPlugin_REM;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_AMO <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_AMO;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_SC <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_SC;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LOAD <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LOAD;
      EU0_ExecutionUnitBase_pipeline_fetch_1_AguPlugin_LR <= EU0_ExecutionUnitBase_pipeline_fetch_0_AguPlugin_LR;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_ECALL <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_ECALL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_EBREAK <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_EBREAK;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_XRET <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_XRET;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_I <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_I;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FENCE_VMA <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FENCE_VMA;
      EU0_ExecutionUnitBase_pipeline_fetch_1_EnvCallPlugin_FLUSH_DATA <= EU0_ExecutionUnitBase_pipeline_fetch_0_EnvCallPlugin_FLUSH_DATA;
      EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_IMM <= EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_IMM;
      EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_MASK <= EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_MASK;
      EU0_ExecutionUnitBase_pipeline_fetch_1_CsrAccessPlugin_CSR_CLEAR <= EU0_ExecutionUnitBase_pipeline_fetch_0_CsrAccessPlugin_CSR_CLEAR;
      EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_REVERT <= EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_REVERT;
      EU0_ExecutionUnitBase_pipeline_fetch_1_SrcStageables_ZERO <= EU0_ExecutionUnitBase_pipeline_fetch_0_SrcStageables_ZERO;
      EU0_ExecutionUnitBase_pipeline_fetch_1_integer_RS2 <= EU0_ExecutionUnitBase_pipeline_fetch_0_integer_RS2;
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_0_ready_output) begin
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_0 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_0;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_1 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_1;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_2 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_2;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_mul_VALUES_3 <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_logic_mul_VALUES_3;
      EU0_ExecutionUnitBase_pipeline_execute_1_DIV_REVERT_RESULT <= EU0_ExecutionUnitBase_pipeline_execute_0_DIV_REVERT_RESULT;
      EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_REM <= EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_REM;
      EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_0_DivPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_1_Frontend_MICRO_OP <= EU0_ExecutionUnitBase_pipeline_execute_0_Frontend_MICRO_OP;
      EU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID <= EU0_ExecutionUnitBase_pipeline_execute_0_ROB_ID;
      EU0_ExecutionUnitBase_pipeline_execute_1_PHYS_RD <= EU0_ExecutionUnitBase_pipeline_execute_0_PHYS_RD;
      EU0_ExecutionUnitBase_pipeline_execute_1_WRITE_RD <= EU0_ExecutionUnitBase_pipeline_execute_0_WRITE_RD;
      EU0_ExecutionUnitBase_pipeline_execute_1_PC <= EU0_ExecutionUnitBase_pipeline_execute_0_PC;
      EU0_ExecutionUnitBase_pipeline_execute_1_CsrAccessPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_0_CsrAccessPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_HIGH <= EU0_ExecutionUnitBase_pipeline_execute_0_MulPlugin_HIGH;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_EBREAK <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_EBREAK;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_ECALL <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_ECALL;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_XRET <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_XRET;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_I <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_I;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FLUSH_DATA <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FLUSH_DATA;
      EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_VMA <= EU0_ExecutionUnitBase_pipeline_execute_0_EnvCallPlugin_FENCE_VMA;
      EU0_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E2 <= EU0_ExecutionUnitBase_pipeline_execute_0_completion_SEL_E2;
    end
    if(EU0_ExecutionUnitBase_pipeline_execute_1_ready_output) begin
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_0_adders_0 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_0;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_logic_steps_0_adders_1 <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_logic_steps_0_adders_1;
      EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_2_DivPlugin_DIV_RESULT <= EU0_ExecutionUnitBase_pipeline_execute_1_DivPlugin_DIV_RESULT;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_2_MulPlugin_HIGH <= EU0_ExecutionUnitBase_pipeline_execute_1_MulPlugin_HIGH;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_EBREAK <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_EBREAK;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_ECALL <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_ECALL;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_XRET <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_XRET;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_I <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_I;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FLUSH_DATA <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FLUSH_DATA;
      EU0_ExecutionUnitBase_pipeline_execute_2_EnvCallPlugin_FENCE_VMA <= EU0_ExecutionUnitBase_pipeline_execute_1_EnvCallPlugin_FENCE_VMA;
      EU0_ExecutionUnitBase_pipeline_execute_2_ROB_ID <= EU0_ExecutionUnitBase_pipeline_execute_1_ROB_ID;
      EU0_ExecutionUnitBase_pipeline_execute_2_PC <= EU0_ExecutionUnitBase_pipeline_execute_1_PC;
      EU0_ExecutionUnitBase_pipeline_execute_2_Frontend_MICRO_OP <= EU0_ExecutionUnitBase_pipeline_execute_1_Frontend_MICRO_OP;
      EU0_ExecutionUnitBase_pipeline_execute_2_CsrAccessPlugin_SEL <= EU0_ExecutionUnitBase_pipeline_execute_1_CsrAccessPlugin_SEL;
      EU0_ExecutionUnitBase_pipeline_execute_2_WRITE_RD <= EU0_ExecutionUnitBase_pipeline_execute_1_WRITE_RD;
      EU0_ExecutionUnitBase_pipeline_execute_2_PHYS_RD <= EU0_ExecutionUnitBase_pipeline_execute_1_PHYS_RD;
      EU0_ExecutionUnitBase_pipeline_execute_2_completion_SEL_E2 <= EU0_ExecutionUnitBase_pipeline_execute_1_completion_SEL_E2;
    end
    DispatchPlugin_logic_pop_0_stagesList_1_OFFSET <= DispatchPlugin_logic_pop_0_stagesList_0_OFFSET;
    DispatchPlugin_logic_pop_0_stagesList_1_UINT <= DispatchPlugin_logic_pop_0_stagesList_0_UINT;
    DispatchPlugin_logic_pop_0_stagesList_1_LATENCY_0 <= DispatchPlugin_logic_pop_0_stagesList_0_LATENCY_0;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_0 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_0;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_1 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_1;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_2 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_2;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_3 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_3;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_4 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_4;
    DispatchPlugin_logic_pop_0_stagesList_1_ALU0_readContext_PHYS_RD_5 <= DispatchPlugin_logic_pop_0_stagesList_0_ALU0_readContext_PHYS_RD_5;
    DispatchPlugin_logic_pop_1_stagesList_1_OFFSET <= DispatchPlugin_logic_pop_1_stagesList_0_OFFSET;
    DispatchPlugin_logic_pop_1_stagesList_1_UINT <= DispatchPlugin_logic_pop_1_stagesList_0_UINT;
    DispatchPlugin_logic_pop_1_stagesList_1_LATENCY_0 <= DispatchPlugin_logic_pop_1_stagesList_0_LATENCY_0;
    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_0 <= DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_0;
    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_1 <= DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_1;
    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_2 <= DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_2;
    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_3 <= DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_3;
    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_4 <= DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_4;
    DispatchPlugin_logic_pop_1_stagesList_1_ALU1_readContext_PHYS_RD_5 <= DispatchPlugin_logic_pop_1_stagesList_0_ALU1_readContext_PHYS_RD_5;
    if(DispatchPlugin_logic_pop_2_stagesList_0_ready_output) begin
      DispatchPlugin_logic_pop_2_stagesList_1_OFFSET <= DispatchPlugin_logic_pop_2_stagesList_0_OFFSET;
      DispatchPlugin_logic_pop_2_stagesList_1_UINT <= DispatchPlugin_logic_pop_2_stagesList_0_UINT;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_0 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_0;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_1 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_1;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_2 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_2;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_3 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_3;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_4 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_4;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_5 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_5;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_6 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_6;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_7 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_7;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_8 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_8;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_9 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_9;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RD_10 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RD_10;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_0 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_0;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_1 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_1;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_2 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_2;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_3 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_3;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_4 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_4;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_5 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_5;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_6 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_6;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_7 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_7;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_8 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_8;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_9 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_9;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_0_10 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_0_10;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_0 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_0;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_1 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_1;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_2 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_2;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_3 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_3;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_4 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_4;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_5 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_5;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_6 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_6;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_7 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_7;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_8 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_8;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_9 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_9;
      DispatchPlugin_logic_pop_2_stagesList_1_EU0_readContext_PHYS_RS_1_10 <= DispatchPlugin_logic_pop_2_stagesList_0_EU0_readContext_PHYS_RS_1_10;
    end
    if(FrontendPlugin_allocated_ready_output) begin
      FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_0 <= FrontendPlugin_allocated_Frontend_DISPATCH_MASK_0;
      FrontendPlugin_dispatch_WRITE_RD_0 <= FrontendPlugin_allocated_WRITE_RD_0;
      FrontendPlugin_dispatch_PHYS_RD_0 <= FrontendPlugin_allocated_PHYS_RD_0;
      FrontendPlugin_dispatch_Frontend_DISPATCH_MASK_1 <= FrontendPlugin_allocated_Frontend_DISPATCH_MASK_1;
      FrontendPlugin_dispatch_WRITE_RD_1 <= FrontendPlugin_allocated_WRITE_RD_1;
      FrontendPlugin_dispatch_PHYS_RD_1 <= FrontendPlugin_allocated_PHYS_RD_1;
      FrontendPlugin_dispatch_BRANCH_ID_0 <= FrontendPlugin_allocated_BRANCH_ID_0;
      FrontendPlugin_dispatch_BRANCH_SEL_0 <= FrontendPlugin_allocated_BRANCH_SEL_0;
      FrontendPlugin_dispatch_BRANCH_ID_1 <= FrontendPlugin_allocated_BRANCH_ID_1;
      FrontendPlugin_dispatch_BRANCH_SEL_1 <= FrontendPlugin_allocated_BRANCH_SEL_1;
      FrontendPlugin_dispatch_ROB_ID <= FrontendPlugin_allocated_ROB_ID;
      FrontendPlugin_dispatch_ARCH_RD_0 <= FrontendPlugin_allocated_ARCH_RD_0;
      FrontendPlugin_dispatch_ARCH_RS_0_0 <= FrontendPlugin_allocated_ARCH_RS_0_0;
      FrontendPlugin_dispatch_READ_RS_0_0 <= FrontendPlugin_allocated_READ_RS_0_0;
      FrontendPlugin_dispatch_PHYS_RS_0_0 <= FrontendPlugin_allocated_PHYS_RS_0_0;
      FrontendPlugin_dispatch_READ_RS_1_0 <= FrontendPlugin_allocated_READ_RS_1_0;
      FrontendPlugin_dispatch_PHYS_RS_1_0 <= FrontendPlugin_allocated_PHYS_RS_1_0;
      FrontendPlugin_dispatch_ARCH_RS_0_1 <= FrontendPlugin_allocated_ARCH_RS_0_1;
      FrontendPlugin_dispatch_READ_RS_0_1 <= FrontendPlugin_allocated_READ_RS_0_1;
      FrontendPlugin_dispatch_PHYS_RS_0_1 <= FrontendPlugin_allocated_PHYS_RS_0_1;
      FrontendPlugin_dispatch_ARCH_RS_1_1 <= FrontendPlugin_allocated_ARCH_RS_1_1;
      FrontendPlugin_dispatch_READ_RS_1_1 <= FrontendPlugin_allocated_READ_RS_1_1;
      FrontendPlugin_dispatch_PHYS_RS_1_1 <= FrontendPlugin_allocated_PHYS_RS_1_1;
      FrontendPlugin_dispatch_BRANCH_HISTORY_0 <= FrontendPlugin_allocated_BRANCH_HISTORY_0;
      FrontendPlugin_dispatch_BRANCH_HISTORY_1 <= FrontendPlugin_allocated_BRANCH_HISTORY_1;
      FrontendPlugin_dispatch_Frontend_MICRO_OP_0 <= FrontendPlugin_allocated_Frontend_MICRO_OP_0;
      FrontendPlugin_dispatch_Frontend_MICRO_OP_1 <= FrontendPlugin_allocated_Frontend_MICRO_OP_1;
      FrontendPlugin_dispatch_LQ_ALLOC_0 <= FrontendPlugin_allocated_LQ_ALLOC_0;
      FrontendPlugin_dispatch_LQ_ALLOC_1 <= FrontendPlugin_allocated_LQ_ALLOC_1;
      FrontendPlugin_dispatch_SQ_ALLOC_0 <= FrontendPlugin_allocated_SQ_ALLOC_0;
      FrontendPlugin_dispatch_SQ_ALLOC_1 <= FrontendPlugin_allocated_SQ_ALLOC_1;
      FrontendPlugin_dispatch_Prediction_IS_BRANCH_0 <= FrontendPlugin_allocated_Prediction_IS_BRANCH_0;
      FrontendPlugin_dispatch_Prediction_IS_BRANCH_1 <= FrontendPlugin_allocated_Prediction_IS_BRANCH_1;
      FrontendPlugin_dispatch_GSHARE_COUNTER_0_0 <= FrontendPlugin_allocated_GSHARE_COUNTER_0_0;
      FrontendPlugin_dispatch_GSHARE_COUNTER_0_1 <= FrontendPlugin_allocated_GSHARE_COUNTER_0_1;
      FrontendPlugin_dispatch_GSHARE_COUNTER_1_0 <= FrontendPlugin_allocated_GSHARE_COUNTER_1_0;
      FrontendPlugin_dispatch_GSHARE_COUNTER_1_1 <= FrontendPlugin_allocated_GSHARE_COUNTER_1_1;
      FrontendPlugin_dispatch_DispatchPlugin_FENCE_OLDER_0 <= FrontendPlugin_allocated_DispatchPlugin_FENCE_OLDER_0;
      FrontendPlugin_dispatch_DispatchPlugin_FENCE_OLDER_1 <= FrontendPlugin_allocated_DispatchPlugin_FENCE_OLDER_1;
      FrontendPlugin_dispatch_DispatchPlugin_FENCE_YOUNGER_0 <= FrontendPlugin_allocated_DispatchPlugin_FENCE_YOUNGER_0;
      FrontendPlugin_dispatch_DispatchPlugin_FENCE_YOUNGER_1 <= FrontendPlugin_allocated_DispatchPlugin_FENCE_YOUNGER_1;
      FrontendPlugin_dispatch_ALU0_ALU1_SEL_0 <= FrontendPlugin_allocated_ALU0_ALU1_SEL_0;
      FrontendPlugin_dispatch_EU0_SEL_0 <= FrontendPlugin_allocated_EU0_SEL_0;
      FrontendPlugin_dispatch_ALU0_ALU1_SEL_1 <= FrontendPlugin_allocated_ALU0_ALU1_SEL_1;
      FrontendPlugin_dispatch_EU0_SEL_1 <= FrontendPlugin_allocated_EU0_SEL_1;
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_0_0 <= FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_0_0;
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_1_0 <= FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_1_0;
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_0_1 <= FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_0_1;
      FrontendPlugin_dispatch_RfDependencyPlugin_setup_SKIP_1_1 <= FrontendPlugin_allocated_RfDependencyPlugin_setup_SKIP_1_1;
    end
    if(FrontendPlugin_decoded_ready_output) begin
      FrontendPlugin_serialized_FETCH_ID_0 <= FrontendPlugin_decoded_FETCH_ID_0;
      FrontendPlugin_serialized_FETCH_ID_1 <= FrontendPlugin_decoded_FETCH_ID_1;
      FrontendPlugin_serialized_READ_RS_0_0 <= FrontendPlugin_decoded_READ_RS_0_0;
      FrontendPlugin_serialized_READ_RS_1_0 <= FrontendPlugin_decoded_READ_RS_1_0;
      FrontendPlugin_serialized_WRITE_RD_0 <= FrontendPlugin_decoded_WRITE_RD_0;
      FrontendPlugin_serialized_ALU0_ALU1_SEL_0 <= FrontendPlugin_decoded_ALU0_ALU1_SEL_0;
      FrontendPlugin_serialized_EU0_SEL_0 <= FrontendPlugin_decoded_EU0_SEL_0;
      FrontendPlugin_serialized_LQ_ALLOC_0 <= FrontendPlugin_decoded_LQ_ALLOC_0;
      FrontendPlugin_serialized_SQ_ALLOC_0 <= FrontendPlugin_decoded_SQ_ALLOC_0;
      FrontendPlugin_serialized_Frontend_DECODED_MASK_0 <= FrontendPlugin_decoded_Frontend_DECODED_MASK_0;
      FrontendPlugin_serialized_Frontend_MICRO_OP_0 <= FrontendPlugin_decoded_Frontend_MICRO_OP_0;
      FrontendPlugin_serialized_ARCH_RD_0 <= FrontendPlugin_decoded_ARCH_RD_0;
      FrontendPlugin_serialized_ARCH_RS_0_0 <= FrontendPlugin_decoded_ARCH_RS_0_0;
      FrontendPlugin_serialized_ARCH_RS_1_0 <= FrontendPlugin_decoded_ARCH_RS_1_0;
      FrontendPlugin_serialized_READ_RS_0_1 <= FrontendPlugin_decoded_READ_RS_0_1;
      FrontendPlugin_serialized_READ_RS_1_1 <= FrontendPlugin_decoded_READ_RS_1_1;
      FrontendPlugin_serialized_WRITE_RD_1 <= FrontendPlugin_decoded_WRITE_RD_1;
      FrontendPlugin_serialized_ALU0_ALU1_SEL_1 <= FrontendPlugin_decoded_ALU0_ALU1_SEL_1;
      FrontendPlugin_serialized_EU0_SEL_1 <= FrontendPlugin_decoded_EU0_SEL_1;
      FrontendPlugin_serialized_LQ_ALLOC_1 <= FrontendPlugin_decoded_LQ_ALLOC_1;
      FrontendPlugin_serialized_SQ_ALLOC_1 <= FrontendPlugin_decoded_SQ_ALLOC_1;
      FrontendPlugin_serialized_Frontend_DECODED_MASK_1 <= FrontendPlugin_decoded_Frontend_DECODED_MASK_1;
      FrontendPlugin_serialized_Frontend_MICRO_OP_1 <= FrontendPlugin_decoded_Frontend_MICRO_OP_1;
      FrontendPlugin_serialized_ARCH_RD_1 <= FrontendPlugin_decoded_ARCH_RD_1;
      FrontendPlugin_serialized_ARCH_RS_0_1 <= FrontendPlugin_decoded_ARCH_RS_0_1;
      FrontendPlugin_serialized_ARCH_RS_1_1 <= FrontendPlugin_decoded_ARCH_RS_1_1;
      FrontendPlugin_serialized_PC_0 <= FrontendPlugin_decoded_PC_0;
      FrontendPlugin_serialized_PC_1 <= FrontendPlugin_decoded_PC_1;
      FrontendPlugin_serialized_OP_ID <= FrontendPlugin_decoded_OP_ID;
      FrontendPlugin_serialized_IS_JALR_0 <= FrontendPlugin_decoded_IS_JALR_0;
      FrontendPlugin_serialized_Prediction_IS_BRANCH_0 <= FrontendPlugin_decoded_Prediction_IS_BRANCH_0;
      FrontendPlugin_serialized_IS_ANY_0 <= FrontendPlugin_decoded_IS_ANY_0;
      FrontendPlugin_serialized_RAS_PUSH_0 <= FrontendPlugin_decoded_RAS_PUSH_0;
      FrontendPlugin_serialized_RAS_POP_0 <= FrontendPlugin_decoded_RAS_POP_0;
      FrontendPlugin_serialized_PC_INC_0 <= FrontendPlugin_decoded_PC_INC_0;
      FrontendPlugin_serialized_PC_TARGET_PRE_RAS_0 <= FrontendPlugin_decoded_PC_TARGET_PRE_RAS_0;
      FrontendPlugin_serialized_BAD_RET_PC_0 <= FrontendPlugin_decoded_BAD_RET_PC_0;
      FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_PC_NEXT_0 <= FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_0;
      FrontendPlugin_serialized_CAN_IMPROVE_0 <= FrontendPlugin_decoded_CAN_IMPROVE_0;
      FrontendPlugin_serialized_BRANCHED_PREDICTION_0 <= FrontendPlugin_decoded_BRANCHED_PREDICTION_0;
      FrontendPlugin_serialized_IS_JALR_1 <= FrontendPlugin_decoded_IS_JALR_1;
      FrontendPlugin_serialized_Prediction_IS_BRANCH_1 <= FrontendPlugin_decoded_Prediction_IS_BRANCH_1;
      FrontendPlugin_serialized_IS_ANY_1 <= FrontendPlugin_decoded_IS_ANY_1;
      FrontendPlugin_serialized_RAS_PUSH_1 <= FrontendPlugin_decoded_RAS_PUSH_1;
      FrontendPlugin_serialized_RAS_POP_1 <= FrontendPlugin_decoded_RAS_POP_1;
      FrontendPlugin_serialized_PC_INC_1 <= FrontendPlugin_decoded_PC_INC_1;
      FrontendPlugin_serialized_PC_TARGET_PRE_RAS_1 <= FrontendPlugin_decoded_PC_TARGET_PRE_RAS_1;
      FrontendPlugin_serialized_BAD_RET_PC_1 <= FrontendPlugin_decoded_BAD_RET_PC_1;
      FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_PC_NEXT_1 <= FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_PC_NEXT_1;
      FrontendPlugin_serialized_CAN_IMPROVE_1 <= FrontendPlugin_decoded_CAN_IMPROVE_1;
      FrontendPlugin_serialized_BRANCHED_PREDICTION_1 <= FrontendPlugin_decoded_BRANCHED_PREDICTION_1;
      FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_0 <= FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_VALID_0;
      FrontendPlugin_serialized_Prediction_ALIGNED_BRANCH_VALID_1 <= FrontendPlugin_decoded_Prediction_ALIGNED_BRANCH_VALID_1;
      FrontendPlugin_serialized_BRANCH_HISTORY_0 <= FrontendPlugin_decoded_BRANCH_HISTORY_0;
      FrontendPlugin_serialized_BRANCH_HISTORY_1 <= FrontendPlugin_decoded_BRANCH_HISTORY_1;
      FrontendPlugin_serialized_GSHARE_COUNTER_0_0 <= FrontendPlugin_decoded_GSHARE_COUNTER_0_0;
      FrontendPlugin_serialized_GSHARE_COUNTER_0_1 <= FrontendPlugin_decoded_GSHARE_COUNTER_0_1;
      FrontendPlugin_serialized_GSHARE_COUNTER_1_0 <= FrontendPlugin_decoded_GSHARE_COUNTER_1_0;
      FrontendPlugin_serialized_GSHARE_COUNTER_1_1 <= FrontendPlugin_decoded_GSHARE_COUNTER_1_1;
    end
    if(FetchPlugin_stages_0_ready_output) begin
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_loaded <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_error <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_error;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_0_address;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_loaded <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_1_loaded;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_error <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_1_error;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_1_address;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_loaded <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_2_loaded;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_error <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_2_error;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_2_address;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_loaded <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_3_loaded;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_error <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_3_error;
      FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address <= FetchPlugin_stages_0_FetchCachePlugin_logic_WAYS_TAGS_3_address;
      FetchPlugin_stages_1_Fetch_FETCH_PC <= FetchPlugin_stages_0_Fetch_FETCH_PC;
      FetchPlugin_stages_1_GSharePlugin_logic_HASH <= FetchPlugin_stages_0_GSharePlugin_logic_HASH;
      FetchPlugin_stages_1_BRANCH_HISTORY <= FetchPlugin_stages_0_BRANCH_HISTORY;
      FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_valid <= FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_valid;
      FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_address <= FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_address;
      FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_data_0 <= FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_data_0;
      FetchPlugin_stages_1_GSharePlugin_logic_BYPASS_payload_data_1 <= FetchPlugin_stages_0_GSharePlugin_logic_BYPASS_payload_data_1;
    end
    if(FetchPlugin_stages_1_ready_output) begin
      FetchPlugin_stages_2_FETCH_ID <= FetchPlugin_stages_1_FETCH_ID;
      FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_0 <= FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_0;
      FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_1 <= FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_1;
      FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_2 <= FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_2;
      FetchPlugin_stages_2_FetchCachePlugin_logic_BANKS_MUXES_3 <= FetchPlugin_stages_1_FetchCachePlugin_logic_BANKS_MUXES_3;
      FetchPlugin_stages_2_Fetch_FETCH_PC <= FetchPlugin_stages_1_Fetch_FETCH_PC;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_loaded <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_loaded;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_error <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_error;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_0_address <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_0_address;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_1_loaded <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_loaded;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_1_error <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_error;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_1_address <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_1_address;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_2_loaded <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_loaded;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_2_error <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_error;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_2_address <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_2_address;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_3_loaded <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_loaded;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_3_error <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_error;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_TAGS_3_address <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_TAGS_3_address;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_0 <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_0;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_1 <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_1;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_2 <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_2;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HITS_3 <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HITS_3;
      FetchPlugin_stages_2_FetchCachePlugin_logic_PLRU_0 <= FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_0;
      FetchPlugin_stages_2_FetchCachePlugin_logic_PLRU_1 <= FetchPlugin_stages_1_FetchCachePlugin_logic_PLRU_1;
      FetchPlugin_stages_2_FetchCachePlugin_logic_WAYS_HIT <= FetchPlugin_stages_1_FetchCachePlugin_logic_WAYS_HIT;
      FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT <= FetchPlugin_stages_1_AlignerPlugin_MASK_FRONT;
      FetchPlugin_stages_2_GSHARE_COUNTER_0 <= FetchPlugin_stages_1_GSHARE_COUNTER_0;
      FetchPlugin_stages_2_GSHARE_COUNTER_1 <= FetchPlugin_stages_1_GSHARE_COUNTER_1;
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID <= FetchPlugin_stages_1_Prediction_WORD_BRANCH_VALID;
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_SLICE <= FetchPlugin_stages_1_Prediction_WORD_BRANCH_SLICE;
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT <= FetchPlugin_stages_1_Prediction_WORD_BRANCH_PC_NEXT;
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID <= FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALID;
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_SLICE <= FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_SLICE;
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE <= FetchPlugin_stages_1_Prediction_BRANCH_HISTORY_PUSH_VALUE;
      FetchPlugin_stages_2_MMU_IO <= FetchPlugin_stages_1_MMU_IO;
      FetchPlugin_stages_2_MMU_TRANSLATED <= FetchPlugin_stages_1_MMU_TRANSLATED;
      FetchPlugin_stages_2_MMU_REDO <= FetchPlugin_stages_1_MMU_REDO;
      FetchPlugin_stages_2_MMU_ALLOW_EXECUTE <= FetchPlugin_stages_1_MMU_ALLOW_EXECUTE;
      FetchPlugin_stages_2_MMU_PAGE_FAULT <= FetchPlugin_stages_1_MMU_PAGE_FAULT;
      FetchPlugin_stages_2_MMU_ACCESS_FAULT <= FetchPlugin_stages_1_MMU_ACCESS_FAULT;
      FetchPlugin_stages_2_Fetch_FETCH_PC_INC <= FetchPlugin_stages_1_Fetch_FETCH_PC_INC;
      FetchPlugin_stages_2_BRANCH_HISTORY <= FetchPlugin_stages_1_BRANCH_HISTORY;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_WORD_s2mBuffer <= FetchPlugin_stages_2_Fetch_WORD;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_FETCH_PC_s2mBuffer <= FetchPlugin_stages_2_Fetch_FETCH_PC;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_WORD_FAULT_s2mBuffer <= FetchPlugin_stages_2_Fetch_WORD_FAULT;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE_s2mBuffer <= FetchPlugin_stages_2_Fetch_WORD_FAULT_PAGE;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_BRANCH_HISTORY_s2mBuffer <= FetchPlugin_stages_2_BRANCH_HISTORY;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_FETCH_ID_s2mBuffer <= FetchPlugin_stages_2_FETCH_ID;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_SLICE_s2mBuffer <= FetchPlugin_stages_2_Prediction_WORD_BRANCH_SLICE;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID_s2mBuffer <= FetchPlugin_stages_2_Prediction_WORD_BRANCH_VALID;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT_s2mBuffer <= FetchPlugin_stages_2_AlignerPlugin_MASK_FRONT;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT_s2mBuffer <= FetchPlugin_stages_2_Prediction_WORD_BRANCH_PC_NEXT;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID_s2mBuffer <= FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALID;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_SLICE_s2mBuffer <= FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_SLICE;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE_s2mBuffer <= FetchPlugin_stages_2_Prediction_BRANCH_HISTORY_PUSH_VALUE;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_GSHARE_COUNTER_s2mBuffer_0 <= FetchPlugin_stages_2_GSHARE_COUNTER_0;
      FetchPlugin_stages_2_GSHARE_COUNTER_s2mBuffer_1 <= FetchPlugin_stages_2_GSHARE_COUNTER_1;
    end
    if(FetchPlugin_stages_2_ready_output) begin
      FetchPlugin_stages_2_Fetch_FETCH_PC_INC_s2mBuffer <= FetchPlugin_stages_2_Fetch_FETCH_PC_INC;
    end
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_enumDef_IDLE : begin
        if(PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
          PerformanceCounterPlugin_logic_fsm_cmd_flusher <= 1'b1;
          PerformanceCounterPlugin_logic_fsm_cmd_address <= PerformanceCounterPlugin_logic_fsm_flusherCmd_payload_address;
        end else begin
          if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
            PerformanceCounterPlugin_logic_fsm_cmd_flusher <= 1'b0;
            PerformanceCounterPlugin_logic_fsm_cmd_address <= PerformanceCounterPlugin_logic_fsm_csrReadCmd_payload_address;
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_LOW : begin
        PerformanceCounterPlugin_logic_fsm_ramReaded[31 : 0] <= PerformanceCounterPlugin_setup_readPort_data;
        PerformanceCounterPlugin_logic_fsm_counterReaded <= _zz_PerformanceCounterPlugin_logic_fsm_counterReaded_11;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CALC : begin
        PerformanceCounterPlugin_logic_fsm_result <= PerformanceCounterPlugin_logic_fsm_calc;
        if(!PerformanceCounterPlugin_logic_fsm_cmd_flusher) begin
          PerformanceCounterPlugin_logic_fsm_resultCsr <= PerformanceCounterPlugin_logic_fsm_calc;
        end
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_READ_HIGH : begin
        PerformanceCounterPlugin_logic_fsm_ramReaded[63 : 32] <= PerformanceCounterPlugin_setup_readPort_data;
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_WRITE_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE : begin
      end
      PerformanceCounterPlugin_logic_fsm_enumDef_CSR_WRITE_COMPLETION : begin
      end
      default : begin
      end
    endcase
    case(PrivilegedPlugin_logic_fsm_stateReg)
      PrivilegedPlugin_logic_fsm_enumDef_IDLE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_SETUP : begin
        if(when_PrivilegedPlugin_l766) begin
          PrivilegedPlugin_logic_fsm_trap_interrupt <= 1'b1;
          PrivilegedPlugin_logic_fsm_trap_code <= PrivilegedPlugin_logic_decoderInterrupt_buffer_code;
          PrivilegedPlugin_logic_fsm_trap_targetPrivilege <= PrivilegedPlugin_logic_decoderInterrupt_buffer_targetPrivilege;
        end else begin
          case(PrivilegedPlugin_logic_reschedule_payload_cause)
            4'b1001 : begin
            end
            4'b1010 : begin
            end
            4'b1000 : begin
            end
            default : begin
              PrivilegedPlugin_logic_fsm_trap_interrupt <= 1'b0;
              PrivilegedPlugin_logic_fsm_trap_code <= PrivilegedPlugin_logic_exception_code;
              PrivilegedPlugin_logic_fsm_trap_targetPrivilege <= PrivilegedPlugin_logic_exception_targetPrivilege;
            end
          endcase
        end
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVAL_WRITE : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_EPC_READ : begin
        PrivilegedPlugin_logic_readed <= PrivilegedPlugin_setup_ramRead_data;
      end
      PrivilegedPlugin_logic_fsm_enumDef_TVEC_READ : begin
        PrivilegedPlugin_logic_readed <= PrivilegedPlugin_setup_ramRead_data;
      end
      PrivilegedPlugin_logic_fsm_enumDef_XRET : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_CALC : begin
        PrivilegedPlugin_logic_readed[31 : 0] <= _zz_PrivilegedPlugin_logic_readed;
      end
      PrivilegedPlugin_logic_fsm_enumDef_FLUSH_JUMP : begin
      end
      PrivilegedPlugin_logic_fsm_enumDef_TRAP : begin
      end
      default : begin
      end
    endcase
    if(Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_cmd_valid) begin
      _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score_3 <= _zz_Lsu2Plugin_logic_aguPush_0_hazardPrediction_read_rsp_score;
    end
    if(Lsu2Plugin_logic_aguPush_0_hitPrediction_read_cmd_valid) begin
      _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter_2 <= _zz_Lsu2Plugin_logic_aguPush_0_hitPrediction_read_rsp_counter;
    end
  end


endmodule

module RamAsyncMwXor_7 (
  input  wire          io_writes_0_valid,
  input  wire [5:0]    io_writes_0_payload_address,
  input  wire [0:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [5:0]    io_writes_1_payload_address,
  input  wire [0:0]    io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [5:0]    io_read_0_cmd_payload,
  output wire [0:0]    io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [5:0]    io_read_1_cmd_payload,
  output wire [0:0]    io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [5:0]    io_read_2_cmd_payload,
  output wire [0:0]    io_read_2_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [0:0]    _zz_ram_0_port1;
  wire       [0:0]    _zz_ram_0_port2;
  wire       [0:0]    _zz_ram_0_port3;
  wire       [0:0]    _zz_ram_0_port4;
  wire       [0:0]    _zz_ram_1_port0;
  wire       [0:0]    _zz_ram_1_port2;
  wire       [0:0]    _zz_ram_1_port3;
  wire       [0:0]    _zz_ram_1_port4;
  wire       [0:0]    writes_0_values_0;
  wire       [0:0]    writes_0_xored;
  wire       [0:0]    writes_1_values_0;
  wire       [0:0]    writes_1_xored;
  wire       [0:0]    reads_0_values_0;
  wire       [0:0]    reads_0_values_1;
  wire       [0:0]    reads_0_xored;
  wire       [0:0]    reads_1_values_0;
  wire       [0:0]    reads_1_values_1;
  wire       [0:0]    reads_1_xored;
  wire       [0:0]    reads_2_values_0;
  wire       [0:0]    reads_2_values_1;
  wire       [0:0]    reads_2_xored;
  (* ram_style = "distributed" *) reg [0:0] ram_0 [0:63];
  (* ram_style = "distributed" *) reg [0:0] ram_1 [0:63];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_0_port3 = ram_0[io_read_1_cmd_payload];
  assign _zz_ram_0_port4 = ram_0[io_read_2_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_1_port3 = ram_1[io_read_1_cmd_payload];
  assign _zz_ram_1_port4 = ram_1[io_read_2_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_xored = (io_writes_0_payload_data ^ writes_0_values_0);
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_xored = (io_writes_1_payload_data ^ writes_1_values_0);
  assign reads_0_values_0 = _zz_ram_0_port2;
  assign reads_0_values_1 = _zz_ram_1_port2;
  assign reads_0_xored = (reads_0_values_0 ^ reads_0_values_1);
  assign io_read_0_rsp = reads_0_xored;
  assign reads_1_values_0 = _zz_ram_0_port3;
  assign reads_1_values_1 = _zz_ram_1_port3;
  assign reads_1_xored = (reads_1_values_0 ^ reads_1_values_1);
  assign io_read_1_rsp = reads_1_xored;
  assign reads_2_values_0 = _zz_ram_0_port4;
  assign reads_2_values_1 = _zz_ram_1_port4;
  assign reads_2_xored = (reads_2_values_0 ^ reads_2_values_1);
  assign io_read_2_rsp = reads_2_xored;

endmodule

module RamAsyncMwMux_2 (
  input  wire          io_writes_0_valid,
  input  wire [3:0]    io_writes_0_payload_address,
  input  wire [28:0]   io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [3:0]    io_writes_1_payload_address,
  input  wire [28:0]   io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [3:0]    io_read_0_cmd_payload,
  output wire [28:0]   io_read_0_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [0:0]    location_io_writes_0_payload_data;
  wire       [0:0]    location_io_writes_1_payload_data;
  wire       [28:0]   _zz_ram_0_port1;
  wire       [28:0]   _zz_ram_1_port1;
  wire       [0:0]    location_io_read_0_rsp;
  reg        [28:0]   _zz_io_read_0_rsp;
  wire       [28:0]   reads_0_reads_0;
  wire       [28:0]   reads_0_reads_1;
  (* ram_style = "distributed" *) reg [28:0] ram_0 [0:15];
  (* ram_style = "distributed" *) reg [28:0] ram_1 [0:15];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= io_writes_0_payload_data;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_read_0_cmd_payload];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= io_writes_1_payload_data;
    end
  end

  assign _zz_ram_1_port1 = ram_1[io_read_0_cmd_payload];
  RamAsyncMwXor_9 location (
    .io_writes_0_valid           (io_writes_0_valid                ), //i
    .io_writes_0_payload_address (io_writes_0_payload_address[3:0] ), //i
    .io_writes_0_payload_data    (location_io_writes_0_payload_data), //i
    .io_writes_1_valid           (io_writes_1_valid                ), //i
    .io_writes_1_payload_address (io_writes_1_payload_address[3:0] ), //i
    .io_writes_1_payload_data    (location_io_writes_1_payload_data), //i
    .io_read_0_cmd_valid         (io_read_0_cmd_valid              ), //i
    .io_read_0_cmd_payload       (io_read_0_cmd_payload[3:0]       ), //i
    .io_read_0_rsp               (location_io_read_0_rsp           ), //o
    .clk                         (clk                              ), //i
    .reset                       (reset                            )  //i
  );
  always @(*) begin
    case(location_io_read_0_rsp)
      1'b0 : _zz_io_read_0_rsp = reads_0_reads_0;
      default : _zz_io_read_0_rsp = reads_0_reads_1;
    endcase
  end

  assign location_io_writes_0_payload_data = 1'b0;
  assign location_io_writes_1_payload_data = 1'b1;
  assign reads_0_reads_0 = _zz_ram_0_port1;
  assign reads_0_reads_1 = _zz_ram_1_port1;
  assign io_read_0_rsp = _zz_io_read_0_rsp;

endmodule

module RamAsyncMwXor_6 (
  input  wire          io_writes_0_valid,
  input  wire [3:0]    io_writes_0_payload_address,
  input  wire [4:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [3:0]    io_writes_1_payload_address,
  input  wire [4:0]    io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [3:0]    io_read_0_cmd_payload,
  output wire [4:0]    io_read_0_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [4:0]    _zz_ram_0_port1;
  wire       [4:0]    _zz_ram_0_port2;
  wire       [4:0]    _zz_ram_1_port0;
  wire       [4:0]    _zz_ram_1_port2;
  wire       [4:0]    writes_0_values_0;
  wire       [4:0]    writes_0_xored;
  wire       [4:0]    writes_1_values_0;
  wire       [4:0]    writes_1_xored;
  wire       [4:0]    reads_0_values_0;
  wire       [4:0]    reads_0_values_1;
  wire       [4:0]    reads_0_xored;
  (* ram_style = "distributed" *) reg [4:0] ram_0 [0:15];
  (* ram_style = "distributed" *) reg [4:0] ram_1 [0:15];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_read_0_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_xored = (io_writes_0_payload_data ^ writes_0_values_0);
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_xored = (io_writes_1_payload_data ^ writes_1_values_0);
  assign reads_0_values_0 = _zz_ram_0_port2;
  assign reads_0_values_1 = _zz_ram_1_port2;
  assign reads_0_xored = (reads_0_values_0 ^ reads_0_values_1);
  assign io_read_0_rsp = reads_0_xored;

endmodule

//RamAsyncMwXor_5 replaced by RamAsyncMwXor_1

//RamAsyncMwXor_4 replaced by RamAsyncMwXor_1

//RamAsyncMwXor_3 replaced by RamAsyncMwXor_10

//RamAsyncMwXor_2 replaced by RamAsyncMwXor_9

module RamAsyncMwXor_1 (
  input  wire          io_writes_0_valid,
  input  wire [3:0]    io_writes_0_payload_address,
  input  wire [0:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [3:0]    io_writes_1_payload_address,
  input  wire [0:0]    io_writes_1_payload_data,
  input  wire          io_writes_2_valid,
  input  wire [3:0]    io_writes_2_payload_address,
  input  wire [0:0]    io_writes_2_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [3:0]    io_read_0_cmd_payload,
  output wire [0:0]    io_read_0_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [0:0]    _zz_ram_0_port1;
  wire       [0:0]    _zz_ram_0_port2;
  wire       [0:0]    _zz_ram_0_port3;
  wire       [0:0]    _zz_ram_1_port0;
  wire       [0:0]    _zz_ram_1_port2;
  wire       [0:0]    _zz_ram_1_port3;
  wire       [0:0]    _zz_ram_2_port0;
  wire       [0:0]    _zz_ram_2_port1;
  wire       [0:0]    _zz_ram_2_port3;
  wire       [0:0]    writes_0_values_0;
  wire       [0:0]    writes_0_values_1;
  wire       [0:0]    writes_0_xored;
  wire       [0:0]    writes_1_values_0;
  wire       [0:0]    writes_1_values_1;
  wire       [0:0]    writes_1_xored;
  wire       [0:0]    writes_2_values_0;
  wire       [0:0]    writes_2_values_1;
  wire       [0:0]    writes_2_xored;
  wire       [0:0]    reads_0_values_0;
  wire       [0:0]    reads_0_values_1;
  wire       [0:0]    reads_0_values_2;
  wire       [0:0]    reads_0_xored;
  (* ram_style = "distributed" *) reg [0:0] ram_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] ram_1 [0:15];
  (* ram_style = "distributed" *) reg [0:0] ram_2 [0:15];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_writes_2_payload_address];
  assign _zz_ram_0_port3 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_writes_2_payload_address];
  assign _zz_ram_1_port3 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_2_port0 = ram_2[io_writes_0_payload_address];
  assign _zz_ram_2_port1 = ram_2[io_writes_1_payload_address];
  always @(posedge clk) begin
    if(io_writes_2_valid) begin
      ram_2[io_writes_2_payload_address] <= writes_2_xored;
    end
  end

  assign _zz_ram_2_port3 = ram_2[io_read_0_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_values_1 = _zz_ram_2_port0;
  assign writes_0_xored = ((io_writes_0_payload_data ^ writes_0_values_0) ^ writes_0_values_1);
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_values_1 = _zz_ram_2_port1;
  assign writes_1_xored = ((io_writes_1_payload_data ^ writes_1_values_0) ^ writes_1_values_1);
  assign writes_2_values_0 = _zz_ram_0_port2;
  assign writes_2_values_1 = _zz_ram_1_port2;
  assign writes_2_xored = ((io_writes_2_payload_data ^ writes_2_values_0) ^ writes_2_values_1);
  assign reads_0_values_0 = _zz_ram_0_port3;
  assign reads_0_values_1 = _zz_ram_1_port3;
  assign reads_0_values_2 = _zz_ram_2_port3;
  assign reads_0_xored = ((reads_0_values_0 ^ reads_0_values_1) ^ reads_0_values_2);
  assign io_read_0_rsp = reads_0_xored;

endmodule

module RamAsyncMwXor (
  input  wire          io_writes_0_valid,
  input  wire [3:0]    io_writes_0_payload_address,
  input  wire [4:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [3:0]    io_writes_1_payload_address,
  input  wire [4:0]    io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [3:0]    io_read_0_cmd_payload,
  output wire [4:0]    io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [3:0]    io_read_1_cmd_payload,
  output wire [4:0]    io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [3:0]    io_read_2_cmd_payload,
  output wire [4:0]    io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [3:0]    io_read_3_cmd_payload,
  output wire [4:0]    io_read_3_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [4:0]    _zz_ram_0_port1;
  wire       [4:0]    _zz_ram_0_port2;
  wire       [4:0]    _zz_ram_0_port3;
  wire       [4:0]    _zz_ram_0_port4;
  wire       [4:0]    _zz_ram_0_port5;
  wire       [4:0]    _zz_ram_1_port0;
  wire       [4:0]    _zz_ram_1_port2;
  wire       [4:0]    _zz_ram_1_port3;
  wire       [4:0]    _zz_ram_1_port4;
  wire       [4:0]    _zz_ram_1_port5;
  wire       [4:0]    writes_0_values_0;
  wire       [4:0]    writes_0_xored;
  wire       [4:0]    writes_1_values_0;
  wire       [4:0]    writes_1_xored;
  wire       [4:0]    reads_0_values_0;
  wire       [4:0]    reads_0_values_1;
  wire       [4:0]    reads_0_xored;
  wire       [4:0]    reads_1_values_0;
  wire       [4:0]    reads_1_values_1;
  wire       [4:0]    reads_1_xored;
  wire       [4:0]    reads_2_values_0;
  wire       [4:0]    reads_2_values_1;
  wire       [4:0]    reads_2_xored;
  wire       [4:0]    reads_3_values_0;
  wire       [4:0]    reads_3_values_1;
  wire       [4:0]    reads_3_xored;
  (* ram_style = "distributed" *) reg [4:0] ram_0 [0:15];
  (* ram_style = "distributed" *) reg [4:0] ram_1 [0:15];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_0_port3 = ram_0[io_read_1_cmd_payload];
  assign _zz_ram_0_port4 = ram_0[io_read_2_cmd_payload];
  assign _zz_ram_0_port5 = ram_0[io_read_3_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_1_port3 = ram_1[io_read_1_cmd_payload];
  assign _zz_ram_1_port4 = ram_1[io_read_2_cmd_payload];
  assign _zz_ram_1_port5 = ram_1[io_read_3_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_xored = (io_writes_0_payload_data ^ writes_0_values_0);
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_xored = (io_writes_1_payload_data ^ writes_1_values_0);
  assign reads_0_values_0 = _zz_ram_0_port2;
  assign reads_0_values_1 = _zz_ram_1_port2;
  assign reads_0_xored = (reads_0_values_0 ^ reads_0_values_1);
  assign io_read_0_rsp = reads_0_xored;
  assign reads_1_values_0 = _zz_ram_0_port3;
  assign reads_1_values_1 = _zz_ram_1_port3;
  assign reads_1_xored = (reads_1_values_0 ^ reads_1_values_1);
  assign io_read_1_rsp = reads_1_xored;
  assign reads_2_values_0 = _zz_ram_0_port4;
  assign reads_2_values_1 = _zz_ram_1_port4;
  assign reads_2_xored = (reads_2_values_0 ^ reads_2_values_1);
  assign io_read_2_rsp = reads_2_xored;
  assign reads_3_values_0 = _zz_ram_0_port5;
  assign reads_3_values_1 = _zz_ram_1_port5;
  assign reads_3_xored = (reads_3_values_0 ^ reads_3_values_1);
  assign io_read_3_rsp = reads_3_xored;

endmodule

module RamAsyncMwMux_1 (
  input  wire          io_writes_0_valid,
  input  wire [3:0]    io_writes_0_payload_address,
  input  wire [64:0]   io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [3:0]    io_writes_1_payload_address,
  input  wire [64:0]   io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [3:0]    io_read_0_cmd_payload,
  output wire [64:0]   io_read_0_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [0:0]    location_io_writes_0_payload_data;
  wire       [0:0]    location_io_writes_1_payload_data;
  wire       [64:0]   _zz_ram_0_port1;
  wire       [64:0]   _zz_ram_1_port1;
  wire       [0:0]    location_io_read_0_rsp;
  reg        [64:0]   _zz_io_read_0_rsp;
  wire       [64:0]   reads_0_reads_0;
  wire       [64:0]   reads_0_reads_1;
  (* ram_style = "distributed" *) reg [64:0] ram_0 [0:15];
  (* ram_style = "distributed" *) reg [64:0] ram_1 [0:15];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= io_writes_0_payload_data;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_read_0_cmd_payload];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= io_writes_1_payload_data;
    end
  end

  assign _zz_ram_1_port1 = ram_1[io_read_0_cmd_payload];
  RamAsyncMwXor_9 location (
    .io_writes_0_valid           (io_writes_0_valid                ), //i
    .io_writes_0_payload_address (io_writes_0_payload_address[3:0] ), //i
    .io_writes_0_payload_data    (location_io_writes_0_payload_data), //i
    .io_writes_1_valid           (io_writes_1_valid                ), //i
    .io_writes_1_payload_address (io_writes_1_payload_address[3:0] ), //i
    .io_writes_1_payload_data    (location_io_writes_1_payload_data), //i
    .io_read_0_cmd_valid         (io_read_0_cmd_valid              ), //i
    .io_read_0_cmd_payload       (io_read_0_cmd_payload[3:0]       ), //i
    .io_read_0_rsp               (location_io_read_0_rsp           ), //o
    .clk                         (clk                              ), //i
    .reset                       (reset                            )  //i
  );
  always @(*) begin
    case(location_io_read_0_rsp)
      1'b0 : _zz_io_read_0_rsp = reads_0_reads_0;
      default : _zz_io_read_0_rsp = reads_0_reads_1;
    endcase
  end

  assign location_io_writes_0_payload_data = 1'b0;
  assign location_io_writes_1_payload_data = 1'b1;
  assign reads_0_reads_0 = _zz_ram_0_port1;
  assign reads_0_reads_1 = _zz_ram_1_port1;
  assign io_read_0_rsp = _zz_io_read_0_rsp;

endmodule

module RamAsyncMwMux (
  input  wire          io_writes_0_valid,
  input  wire [3:0]    io_writes_0_payload_address,
  input  wire [32:0]   io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [3:0]    io_writes_1_payload_address,
  input  wire [32:0]   io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [3:0]    io_read_0_cmd_payload,
  output wire [32:0]   io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [3:0]    io_read_1_cmd_payload,
  output wire [32:0]   io_read_1_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [0:0]    location_io_writes_0_payload_data;
  wire       [0:0]    location_io_writes_1_payload_data;
  wire       [32:0]   _zz_ram_0_port1;
  wire       [32:0]   _zz_ram_0_port2;
  wire       [32:0]   _zz_ram_1_port1;
  wire       [32:0]   _zz_ram_1_port2;
  wire       [0:0]    location_io_read_0_rsp;
  wire       [0:0]    location_io_read_1_rsp;
  reg        [32:0]   _zz_io_read_0_rsp;
  reg        [32:0]   _zz_io_read_1_rsp;
  wire       [32:0]   reads_0_reads_0;
  wire       [32:0]   reads_0_reads_1;
  wire       [32:0]   reads_1_reads_0;
  wire       [32:0]   reads_1_reads_1;
  (* ram_style = "distributed" *) reg [32:0] ram_0 [0:15];
  (* ram_style = "distributed" *) reg [32:0] ram_1 [0:15];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= io_writes_0_payload_data;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_0_port2 = ram_0[io_read_1_cmd_payload];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= io_writes_1_payload_data;
    end
  end

  assign _zz_ram_1_port1 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_1_port2 = ram_1[io_read_1_cmd_payload];
  RamAsyncMwXor_10 location (
    .io_writes_0_valid           (io_writes_0_valid                ), //i
    .io_writes_0_payload_address (io_writes_0_payload_address[3:0] ), //i
    .io_writes_0_payload_data    (location_io_writes_0_payload_data), //i
    .io_writes_1_valid           (io_writes_1_valid                ), //i
    .io_writes_1_payload_address (io_writes_1_payload_address[3:0] ), //i
    .io_writes_1_payload_data    (location_io_writes_1_payload_data), //i
    .io_read_0_cmd_valid         (io_read_0_cmd_valid              ), //i
    .io_read_0_cmd_payload       (io_read_0_cmd_payload[3:0]       ), //i
    .io_read_0_rsp               (location_io_read_0_rsp           ), //o
    .io_read_1_cmd_valid         (io_read_1_cmd_valid              ), //i
    .io_read_1_cmd_payload       (io_read_1_cmd_payload[3:0]       ), //i
    .io_read_1_rsp               (location_io_read_1_rsp           ), //o
    .clk                         (clk                              ), //i
    .reset                       (reset                            )  //i
  );
  always @(*) begin
    case(location_io_read_0_rsp)
      1'b0 : _zz_io_read_0_rsp = reads_0_reads_0;
      default : _zz_io_read_0_rsp = reads_0_reads_1;
    endcase
  end

  always @(*) begin
    case(location_io_read_1_rsp)
      1'b0 : _zz_io_read_1_rsp = reads_1_reads_0;
      default : _zz_io_read_1_rsp = reads_1_reads_1;
    endcase
  end

  assign location_io_writes_0_payload_data = 1'b0;
  assign location_io_writes_1_payload_data = 1'b1;
  assign reads_0_reads_0 = _zz_ram_0_port1;
  assign reads_0_reads_1 = _zz_ram_1_port1;
  assign io_read_0_rsp = _zz_io_read_0_rsp;
  assign reads_1_reads_0 = _zz_ram_0_port2;
  assign reads_1_reads_1 = _zz_ram_1_port2;
  assign io_read_1_rsp = _zz_io_read_1_rsp;

endmodule

module DependencyStorage (
  input  wire          io_writes_0_valid,
  input  wire [5:0]    io_writes_0_payload_physical,
  input  wire [5:0]    io_writes_0_payload_robId,
  input  wire          io_writes_1_valid,
  input  wire [5:0]    io_writes_1_payload_physical,
  input  wire [5:0]    io_writes_1_payload_robId,
  input  wire          io_commits_0_valid,
  input  wire [5:0]    io_commits_0_payload_physical,
  input  wire          io_commits_1_valid,
  input  wire [5:0]    io_commits_1_payload_physical,
  input  wire          io_commits_2_valid,
  input  wire [5:0]    io_commits_2_payload_physical,
  input  wire          io_commits_3_valid,
  input  wire [5:0]    io_commits_3_payload_physical,
  input  wire          io_commits_4_valid,
  input  wire [5:0]    io_commits_4_payload_physical,
  input  wire          io_commits_5_valid,
  input  wire [5:0]    io_commits_5_payload_physical,
  input  wire          io_reads_0_cmd_valid,
  input  wire [5:0]    io_reads_0_cmd_payload,
  output wire          io_reads_0_rsp_valid,
  output wire          io_reads_0_rsp_payload_enable,
  output wire [5:0]    io_reads_0_rsp_payload_rob,
  input  wire          io_reads_1_cmd_valid,
  input  wire [5:0]    io_reads_1_cmd_payload,
  output wire          io_reads_1_rsp_valid,
  output wire          io_reads_1_rsp_payload_enable,
  output wire [5:0]    io_reads_1_rsp_payload_rob,
  input  wire          io_reads_2_cmd_valid,
  input  wire [5:0]    io_reads_2_cmd_payload,
  output wire          io_reads_2_rsp_valid,
  output wire          io_reads_2_rsp_payload_enable,
  output wire [5:0]    io_reads_2_rsp_payload_rob,
  input  wire          io_reads_3_cmd_valid,
  input  wire [5:0]    io_reads_3_cmd_payload,
  output wire          io_reads_3_rsp_valid,
  output wire          io_reads_3_rsp_payload_enable,
  output wire [5:0]    io_reads_3_rsp_payload_rob,
  input  wire          clk,
  input  wire          reset
);

  wire       [5:0]    translation_physToRob_io_writes_0_payload_data;
  wire       [5:0]    translation_physToRob_io_writes_1_payload_data;
  wire                translation_physToRob_io_read_0_cmd_valid;
  wire                translation_physToRob_io_read_1_cmd_valid;
  wire                translation_physToRob_io_read_2_cmd_valid;
  wire                translation_physToRob_io_read_3_cmd_valid;
  wire       [0:0]    status_busy_io_writes_0_payload_data;
  wire       [0:0]    status_busy_io_writes_1_payload_data;
  wire       [0:0]    status_busy_io_writes_2_payload_data;
  wire       [0:0]    status_busy_io_writes_3_payload_data;
  wire       [0:0]    status_busy_io_writes_4_payload_data;
  wire       [0:0]    status_busy_io_writes_5_payload_data;
  wire       [0:0]    status_busy_io_writes_6_payload_data;
  wire       [0:0]    status_busy_io_writes_7_payload_data;
  wire                status_busy_io_read_0_cmd_valid;
  wire                status_busy_io_read_1_cmd_valid;
  wire                status_busy_io_read_2_cmd_valid;
  wire                status_busy_io_read_3_cmd_valid;
  wire       [5:0]    translation_physToRob_io_read_0_rsp;
  wire       [5:0]    translation_physToRob_io_read_1_rsp;
  wire       [5:0]    translation_physToRob_io_read_2_rsp;
  wire       [5:0]    translation_physToRob_io_read_3_rsp;
  wire       [0:0]    status_busy_io_read_0_rsp;
  wire       [0:0]    status_busy_io_read_1_rsp;
  wire       [0:0]    status_busy_io_read_2_rsp;
  wire       [0:0]    status_busy_io_read_3_rsp;
  wire       [5:0]    read_0_robId;
  wire                read_0_enabled;
  wire       [5:0]    read_1_robId;
  wire                read_1_enabled;
  wire       [5:0]    read_2_robId;
  wire                read_2_enabled;
  wire       [5:0]    read_3_robId;
  wire                read_3_enabled;

  RamAsyncMwXor_11 translation_physToRob (
    .io_writes_0_valid           (io_writes_0_valid                                  ), //i
    .io_writes_0_payload_address (io_writes_0_payload_physical[5:0]                  ), //i
    .io_writes_0_payload_data    (translation_physToRob_io_writes_0_payload_data[5:0]), //i
    .io_writes_1_valid           (io_writes_1_valid                                  ), //i
    .io_writes_1_payload_address (io_writes_1_payload_physical[5:0]                  ), //i
    .io_writes_1_payload_data    (translation_physToRob_io_writes_1_payload_data[5:0]), //i
    .io_read_0_cmd_valid         (translation_physToRob_io_read_0_cmd_valid          ), //i
    .io_read_0_cmd_payload       (io_reads_0_cmd_payload[5:0]                        ), //i
    .io_read_0_rsp               (translation_physToRob_io_read_0_rsp[5:0]           ), //o
    .io_read_1_cmd_valid         (translation_physToRob_io_read_1_cmd_valid          ), //i
    .io_read_1_cmd_payload       (io_reads_1_cmd_payload[5:0]                        ), //i
    .io_read_1_rsp               (translation_physToRob_io_read_1_rsp[5:0]           ), //o
    .io_read_2_cmd_valid         (translation_physToRob_io_read_2_cmd_valid          ), //i
    .io_read_2_cmd_payload       (io_reads_2_cmd_payload[5:0]                        ), //i
    .io_read_2_rsp               (translation_physToRob_io_read_2_rsp[5:0]           ), //o
    .io_read_3_cmd_valid         (translation_physToRob_io_read_3_cmd_valid          ), //i
    .io_read_3_cmd_payload       (io_reads_3_cmd_payload[5:0]                        ), //i
    .io_read_3_rsp               (translation_physToRob_io_read_3_rsp[5:0]           ), //o
    .clk                         (clk                                                ), //i
    .reset                       (reset                                              )  //i
  );
  RamAsyncMwXor_12 status_busy (
    .io_writes_0_valid           (io_writes_0_valid                   ), //i
    .io_writes_0_payload_address (io_writes_0_payload_physical[5:0]   ), //i
    .io_writes_0_payload_data    (status_busy_io_writes_0_payload_data), //i
    .io_writes_1_valid           (io_writes_1_valid                   ), //i
    .io_writes_1_payload_address (io_writes_1_payload_physical[5:0]   ), //i
    .io_writes_1_payload_data    (status_busy_io_writes_1_payload_data), //i
    .io_writes_2_valid           (io_commits_0_valid                  ), //i
    .io_writes_2_payload_address (io_commits_0_payload_physical[5:0]  ), //i
    .io_writes_2_payload_data    (status_busy_io_writes_2_payload_data), //i
    .io_writes_3_valid           (io_commits_1_valid                  ), //i
    .io_writes_3_payload_address (io_commits_1_payload_physical[5:0]  ), //i
    .io_writes_3_payload_data    (status_busy_io_writes_3_payload_data), //i
    .io_writes_4_valid           (io_commits_2_valid                  ), //i
    .io_writes_4_payload_address (io_commits_2_payload_physical[5:0]  ), //i
    .io_writes_4_payload_data    (status_busy_io_writes_4_payload_data), //i
    .io_writes_5_valid           (io_commits_3_valid                  ), //i
    .io_writes_5_payload_address (io_commits_3_payload_physical[5:0]  ), //i
    .io_writes_5_payload_data    (status_busy_io_writes_5_payload_data), //i
    .io_writes_6_valid           (io_commits_4_valid                  ), //i
    .io_writes_6_payload_address (io_commits_4_payload_physical[5:0]  ), //i
    .io_writes_6_payload_data    (status_busy_io_writes_6_payload_data), //i
    .io_writes_7_valid           (io_commits_5_valid                  ), //i
    .io_writes_7_payload_address (io_commits_5_payload_physical[5:0]  ), //i
    .io_writes_7_payload_data    (status_busy_io_writes_7_payload_data), //i
    .io_read_0_cmd_valid         (status_busy_io_read_0_cmd_valid     ), //i
    .io_read_0_cmd_payload       (io_reads_0_cmd_payload[5:0]         ), //i
    .io_read_0_rsp               (status_busy_io_read_0_rsp           ), //o
    .io_read_1_cmd_valid         (status_busy_io_read_1_cmd_valid     ), //i
    .io_read_1_cmd_payload       (io_reads_1_cmd_payload[5:0]         ), //i
    .io_read_1_rsp               (status_busy_io_read_1_rsp           ), //o
    .io_read_2_cmd_valid         (status_busy_io_read_2_cmd_valid     ), //i
    .io_read_2_cmd_payload       (io_reads_2_cmd_payload[5:0]         ), //i
    .io_read_2_rsp               (status_busy_io_read_2_rsp           ), //o
    .io_read_3_cmd_valid         (status_busy_io_read_3_cmd_valid     ), //i
    .io_read_3_cmd_payload       (io_reads_3_cmd_payload[5:0]         ), //i
    .io_read_3_rsp               (status_busy_io_read_3_rsp           ), //o
    .clk                         (clk                                 ), //i
    .reset                       (reset                               )  //i
  );
  assign read_0_robId = translation_physToRob_io_read_0_rsp;
  assign read_0_enabled = status_busy_io_read_0_rsp[0];
  assign io_reads_0_rsp_valid = io_reads_0_cmd_valid;
  assign io_reads_0_rsp_payload_enable = read_0_enabled;
  assign io_reads_0_rsp_payload_rob = read_0_robId;
  assign read_1_robId = translation_physToRob_io_read_1_rsp;
  assign read_1_enabled = status_busy_io_read_1_rsp[0];
  assign io_reads_1_rsp_valid = io_reads_1_cmd_valid;
  assign io_reads_1_rsp_payload_enable = read_1_enabled;
  assign io_reads_1_rsp_payload_rob = read_1_robId;
  assign read_2_robId = translation_physToRob_io_read_2_rsp;
  assign read_2_enabled = status_busy_io_read_2_rsp[0];
  assign io_reads_2_rsp_valid = io_reads_2_cmd_valid;
  assign io_reads_2_rsp_payload_enable = read_2_enabled;
  assign io_reads_2_rsp_payload_rob = read_2_robId;
  assign read_3_robId = translation_physToRob_io_read_3_rsp;
  assign read_3_enabled = status_busy_io_read_3_rsp[0];
  assign io_reads_3_rsp_valid = io_reads_3_cmd_valid;
  assign io_reads_3_rsp_payload_enable = read_3_enabled;
  assign io_reads_3_rsp_payload_rob = read_3_robId;
  assign translation_physToRob_io_writes_0_payload_data = io_writes_0_payload_robId;
  assign translation_physToRob_io_writes_1_payload_data = io_writes_1_payload_robId;
  assign translation_physToRob_io_read_0_cmd_valid = 1'b1;
  assign translation_physToRob_io_read_1_cmd_valid = 1'b1;
  assign translation_physToRob_io_read_2_cmd_valid = 1'b1;
  assign translation_physToRob_io_read_3_cmd_valid = 1'b1;
  assign status_busy_io_writes_0_payload_data = 1'b1;
  assign status_busy_io_writes_1_payload_data = 1'b1;
  assign status_busy_io_writes_2_payload_data = 1'b0;
  assign status_busy_io_writes_3_payload_data = 1'b0;
  assign status_busy_io_writes_4_payload_data = 1'b0;
  assign status_busy_io_writes_5_payload_data = 1'b0;
  assign status_busy_io_writes_6_payload_data = 1'b0;
  assign status_busy_io_writes_7_payload_data = 1'b0;
  assign status_busy_io_read_0_cmd_valid = 1'b1;
  assign status_busy_io_read_1_cmd_valid = 1'b1;
  assign status_busy_io_read_2_cmd_valid = 1'b1;
  assign status_busy_io_read_3_cmd_valid = 1'b1;

endmodule

module RegFileAsync (
  input  wire          io_writes_0_valid,
  input  wire [5:0]    io_writes_0_address,
  input  wire [31:0]   io_writes_0_data,
  input  wire [5:0]    io_writes_0_robId,
  input  wire          io_writes_1_valid,
  input  wire [5:0]    io_writes_1_address,
  input  wire [31:0]   io_writes_1_data,
  input  wire [5:0]    io_writes_1_robId,
  input  wire          io_writes_2_valid,
  input  wire [5:0]    io_writes_2_address,
  input  wire [31:0]   io_writes_2_data,
  input  wire [5:0]    io_writes_2_robId,
  input  wire          io_writes_3_valid,
  input  wire [5:0]    io_writes_3_address,
  input  wire [31:0]   io_writes_3_data,
  input  wire [5:0]    io_writes_3_robId,
  input  wire          io_reads_0_valid,
  input  wire [5:0]    io_reads_0_address,
  output wire [31:0]   io_reads_0_data,
  input  wire          io_reads_1_valid,
  input  wire [5:0]    io_reads_1_address,
  output wire [31:0]   io_reads_1_data,
  input  wire          io_reads_2_valid,
  input  wire [5:0]    io_reads_2_address,
  output wire [31:0]   io_reads_2_data,
  input  wire          io_reads_3_valid,
  input  wire [5:0]    io_reads_3_address,
  output wire [31:0]   io_reads_3_data,
  input  wire          io_reads_4_valid,
  input  wire [5:0]    io_reads_4_address,
  output wire [31:0]   io_reads_4_data,
  input  wire          io_reads_5_valid,
  input  wire [5:0]    io_reads_5_address,
  output wire [31:0]   io_reads_5_data,
  input  wire          clk,
  input  wire          reset
);

  wire                banks_0_ram_io_read_0_cmd_valid;
  wire                banks_0_ram_io_read_1_cmd_valid;
  wire                banks_0_ram_io_read_2_cmd_valid;
  wire                banks_0_ram_io_read_3_cmd_valid;
  wire                banks_0_ram_io_read_4_cmd_valid;
  wire                banks_0_ram_io_read_5_cmd_valid;
  wire       [31:0]   banks_0_ram_io_read_0_rsp;
  wire       [31:0]   banks_0_ram_io_read_1_rsp;
  wire       [31:0]   banks_0_ram_io_read_2_rsp;
  wire       [31:0]   banks_0_ram_io_read_3_rsp;
  wire       [31:0]   banks_0_ram_io_read_4_rsp;
  wire       [31:0]   banks_0_ram_io_read_5_rsp;
  reg                 _zz_io_writes_3_valid;
  reg                 _zz_io_writes_2_valid;
  reg                 _zz_io_writes_1_valid;
  reg                 _zz_io_writes_0_valid;
  wire                banks_0_writePort_0_valid;
  wire       [5:0]    banks_0_writePort_0_payload_address;
  wire       [31:0]   banks_0_writePort_0_payload_data;
  reg                 banks_0_writePort_1_valid;
  reg        [5:0]    banks_0_writePort_1_payload_address;
  reg        [31:0]   banks_0_writePort_1_payload_data;
  wire                banks_0_writePort_2_valid;
  wire       [5:0]    banks_0_writePort_2_payload_address;
  wire       [31:0]   banks_0_writePort_2_payload_data;
  wire                banks_0_writePort_3_valid;
  wire       [5:0]    banks_0_writePort_3_payload_address;
  wire       [31:0]   banks_0_writePort_3_payload_data;
  wire       [5:0]    banks_0_readPort_0_address;
  wire       [31:0]   banks_0_readPort_0_data;
  wire       [5:0]    banks_0_readPort_1_address;
  wire       [31:0]   banks_0_readPort_1_data;
  wire       [5:0]    banks_0_readPort_2_address;
  wire       [31:0]   banks_0_readPort_2_data;
  wire       [5:0]    banks_0_readPort_3_address;
  wire       [31:0]   banks_0_readPort_3_data;
  wire       [5:0]    banks_0_readPort_4_address;
  wire       [31:0]   banks_0_readPort_4_data;
  wire       [5:0]    banks_0_readPort_5_address;
  wire       [31:0]   banks_0_readPort_5_data;
  reg                 initHead_booted;
  wire                when_RegFilePlugin_l77;

  RamAsyncMwMux_3 banks_0_ram (
    .io_writes_0_valid           (_zz_io_writes_0_valid                   ), //i
    .io_writes_0_payload_address (banks_0_writePort_0_payload_address[5:0]), //i
    .io_writes_0_payload_data    (banks_0_writePort_0_payload_data[31:0]  ), //i
    .io_writes_1_valid           (_zz_io_writes_1_valid                   ), //i
    .io_writes_1_payload_address (banks_0_writePort_1_payload_address[5:0]), //i
    .io_writes_1_payload_data    (banks_0_writePort_1_payload_data[31:0]  ), //i
    .io_writes_2_valid           (_zz_io_writes_2_valid                   ), //i
    .io_writes_2_payload_address (banks_0_writePort_2_payload_address[5:0]), //i
    .io_writes_2_payload_data    (banks_0_writePort_2_payload_data[31:0]  ), //i
    .io_writes_3_valid           (_zz_io_writes_3_valid                   ), //i
    .io_writes_3_payload_address (banks_0_writePort_3_payload_address[5:0]), //i
    .io_writes_3_payload_data    (banks_0_writePort_3_payload_data[31:0]  ), //i
    .io_read_0_cmd_valid         (banks_0_ram_io_read_0_cmd_valid         ), //i
    .io_read_0_cmd_payload       (banks_0_readPort_0_address[5:0]         ), //i
    .io_read_0_rsp               (banks_0_ram_io_read_0_rsp[31:0]         ), //o
    .io_read_1_cmd_valid         (banks_0_ram_io_read_1_cmd_valid         ), //i
    .io_read_1_cmd_payload       (banks_0_readPort_1_address[5:0]         ), //i
    .io_read_1_rsp               (banks_0_ram_io_read_1_rsp[31:0]         ), //o
    .io_read_2_cmd_valid         (banks_0_ram_io_read_2_cmd_valid         ), //i
    .io_read_2_cmd_payload       (banks_0_readPort_2_address[5:0]         ), //i
    .io_read_2_rsp               (banks_0_ram_io_read_2_rsp[31:0]         ), //o
    .io_read_3_cmd_valid         (banks_0_ram_io_read_3_cmd_valid         ), //i
    .io_read_3_cmd_payload       (banks_0_readPort_3_address[5:0]         ), //i
    .io_read_3_rsp               (banks_0_ram_io_read_3_rsp[31:0]         ), //o
    .io_read_4_cmd_valid         (banks_0_ram_io_read_4_cmd_valid         ), //i
    .io_read_4_cmd_payload       (banks_0_readPort_4_address[5:0]         ), //i
    .io_read_4_rsp               (banks_0_ram_io_read_4_rsp[31:0]         ), //o
    .io_read_5_cmd_valid         (banks_0_ram_io_read_5_cmd_valid         ), //i
    .io_read_5_cmd_payload       (banks_0_readPort_5_address[5:0]         ), //i
    .io_read_5_rsp               (banks_0_ram_io_read_5_rsp[31:0]         ), //o
    .clk                         (clk                                     ), //i
    .reset                       (reset                                   )  //i
  );
  always @(*) begin
    _zz_io_writes_3_valid = 1'b0;
    if(banks_0_writePort_3_valid) begin
      _zz_io_writes_3_valid = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_writes_2_valid = 1'b0;
    if(banks_0_writePort_2_valid) begin
      _zz_io_writes_2_valid = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_writes_1_valid = 1'b0;
    if(banks_0_writePort_1_valid) begin
      _zz_io_writes_1_valid = 1'b1;
    end
  end

  always @(*) begin
    _zz_io_writes_0_valid = 1'b0;
    if(banks_0_writePort_0_valid) begin
      _zz_io_writes_0_valid = 1'b1;
    end
  end

  assign banks_0_readPort_0_data = banks_0_ram_io_read_0_rsp;
  assign banks_0_readPort_1_data = banks_0_ram_io_read_1_rsp;
  assign banks_0_readPort_2_data = banks_0_ram_io_read_2_rsp;
  assign banks_0_readPort_3_data = banks_0_ram_io_read_3_rsp;
  assign banks_0_readPort_4_data = banks_0_ram_io_read_4_rsp;
  assign banks_0_readPort_5_data = banks_0_ram_io_read_5_rsp;
  assign banks_0_writePort_0_valid = (io_writes_0_valid && 1'b1);
  assign banks_0_writePort_0_payload_address = io_writes_0_address;
  assign banks_0_writePort_0_payload_data = io_writes_0_data;
  always @(*) begin
    banks_0_writePort_1_valid = (io_writes_1_valid && 1'b1);
    if(when_RegFilePlugin_l77) begin
      banks_0_writePort_1_valid = 1'b1;
    end
  end

  always @(*) begin
    banks_0_writePort_1_payload_address = io_writes_1_address;
    if(when_RegFilePlugin_l77) begin
      banks_0_writePort_1_payload_address = 6'h00;
    end
  end

  always @(*) begin
    banks_0_writePort_1_payload_data = io_writes_1_data;
    if(when_RegFilePlugin_l77) begin
      banks_0_writePort_1_payload_data = 32'h00000000;
    end
  end

  assign banks_0_writePort_2_valid = (io_writes_2_valid && 1'b1);
  assign banks_0_writePort_2_payload_address = io_writes_2_address;
  assign banks_0_writePort_2_payload_data = io_writes_2_data;
  assign banks_0_writePort_3_valid = (io_writes_3_valid && 1'b1);
  assign banks_0_writePort_3_payload_address = io_writes_3_address;
  assign banks_0_writePort_3_payload_data = io_writes_3_data;
  assign banks_0_readPort_0_address = io_reads_0_address;
  assign io_reads_0_data = banks_0_readPort_0_data;
  assign banks_0_readPort_1_address = io_reads_1_address;
  assign io_reads_1_data = banks_0_readPort_1_data;
  assign banks_0_readPort_2_address = io_reads_2_address;
  assign io_reads_2_data = banks_0_readPort_2_data;
  assign banks_0_readPort_3_address = io_reads_3_address;
  assign io_reads_3_data = banks_0_readPort_3_data;
  assign banks_0_readPort_4_address = io_reads_4_address;
  assign io_reads_4_data = banks_0_readPort_4_data;
  assign banks_0_readPort_5_address = io_reads_5_address;
  assign io_reads_5_data = banks_0_readPort_5_data;
  assign when_RegFilePlugin_l77 = (! initHead_booted);
  assign banks_0_ram_io_read_0_cmd_valid = 1'b1;
  assign banks_0_ram_io_read_1_cmd_valid = 1'b1;
  assign banks_0_ram_io_read_2_cmd_valid = 1'b1;
  assign banks_0_ram_io_read_3_cmd_valid = 1'b1;
  assign banks_0_ram_io_read_4_cmd_valid = 1'b1;
  assign banks_0_ram_io_read_5_cmd_valid = 1'b1;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      initHead_booted <= 1'b0;
    end else begin
      initHead_booted <= 1'b1;
    end
  end


endmodule

module IssueQueue (
  input  wire          io_clear,
  (* keep , syn_keep *) input  wire [31:0]   io_events /* synthesis syn_keep = 1 */ ,
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_slots_0_event,
  input  wire [1:0]    io_push_payload_slots_0_sel,
  input  wire [0:0]    io_push_payload_slots_0_context_staticWake,
  input  wire [5:0]    io_push_payload_slots_0_context_physRd,
  input  wire [5:0]    io_push_payload_slots_0_context_robId,
  input  wire [5:0]    io_push_payload_slots_0_context_euCtx_0,
  input  wire [5:0]    io_push_payload_slots_0_context_euCtx_1,
  input  wire [31:0]   io_push_payload_slots_1_event,
  input  wire [1:0]    io_push_payload_slots_1_sel,
  input  wire [0:0]    io_push_payload_slots_1_context_staticWake,
  input  wire [5:0]    io_push_payload_slots_1_context_physRd,
  input  wire [5:0]    io_push_payload_slots_1_context_robId,
  input  wire [5:0]    io_push_payload_slots_1_context_euCtx_0,
  input  wire [5:0]    io_push_payload_slots_1_context_euCtx_1,
  output wire          io_schedules_0_valid,
  input  wire          io_schedules_0_ready,
  output wire [15:0]   io_schedules_0_payload_event,
  output wire          io_schedules_1_valid,
  input  wire          io_schedules_1_ready,
  output wire [15:0]   io_schedules_1_payload_event,
  output wire          io_schedules_2_valid,
  input  wire          io_schedules_2_ready,
  output wire [31:0]   io_schedules_2_payload_event,
  output wire [0:0]    io_contexts_0_staticWake,
  output wire [5:0]    io_contexts_0_physRd,
  output wire [5:0]    io_contexts_0_robId,
  output wire [5:0]    io_contexts_0_euCtx_0,
  output wire [5:0]    io_contexts_0_euCtx_1,
  output wire [0:0]    io_contexts_1_staticWake,
  output wire [5:0]    io_contexts_1_physRd,
  output wire [5:0]    io_contexts_1_robId,
  output wire [5:0]    io_contexts_1_euCtx_0,
  output wire [5:0]    io_contexts_1_euCtx_1,
  output wire [0:0]    io_contexts_2_staticWake,
  output wire [5:0]    io_contexts_2_physRd,
  output wire [5:0]    io_contexts_2_robId,
  output wire [5:0]    io_contexts_2_euCtx_0,
  output wire [5:0]    io_contexts_2_euCtx_1,
  output wire [0:0]    io_contexts_3_staticWake,
  output wire [5:0]    io_contexts_3_physRd,
  output wire [5:0]    io_contexts_3_robId,
  output wire [5:0]    io_contexts_3_euCtx_0,
  output wire [5:0]    io_contexts_3_euCtx_1,
  output wire [0:0]    io_contexts_4_staticWake,
  output wire [5:0]    io_contexts_4_physRd,
  output wire [5:0]    io_contexts_4_robId,
  output wire [5:0]    io_contexts_4_euCtx_0,
  output wire [5:0]    io_contexts_4_euCtx_1,
  output wire [0:0]    io_contexts_5_staticWake,
  output wire [5:0]    io_contexts_5_physRd,
  output wire [5:0]    io_contexts_5_robId,
  output wire [5:0]    io_contexts_5_euCtx_0,
  output wire [5:0]    io_contexts_5_euCtx_1,
  output wire [0:0]    io_contexts_6_staticWake,
  output wire [5:0]    io_contexts_6_physRd,
  output wire [5:0]    io_contexts_6_robId,
  output wire [5:0]    io_contexts_6_euCtx_0,
  output wire [5:0]    io_contexts_6_euCtx_1,
  output wire [0:0]    io_contexts_7_staticWake,
  output wire [5:0]    io_contexts_7_physRd,
  output wire [5:0]    io_contexts_7_robId,
  output wire [5:0]    io_contexts_7_euCtx_0,
  output wire [5:0]    io_contexts_7_euCtx_1,
  output wire [0:0]    io_contexts_8_staticWake,
  output wire [5:0]    io_contexts_8_physRd,
  output wire [5:0]    io_contexts_8_robId,
  output wire [5:0]    io_contexts_8_euCtx_0,
  output wire [5:0]    io_contexts_8_euCtx_1,
  output wire [0:0]    io_contexts_9_staticWake,
  output wire [5:0]    io_contexts_9_physRd,
  output wire [5:0]    io_contexts_9_robId,
  output wire [5:0]    io_contexts_9_euCtx_0,
  output wire [5:0]    io_contexts_9_euCtx_1,
  output wire [0:0]    io_contexts_10_staticWake,
  output wire [5:0]    io_contexts_10_physRd,
  output wire [5:0]    io_contexts_10_robId,
  output wire [5:0]    io_contexts_10_euCtx_0,
  output wire [5:0]    io_contexts_10_euCtx_1,
  output wire [0:0]    io_contexts_11_staticWake,
  output wire [5:0]    io_contexts_11_physRd,
  output wire [5:0]    io_contexts_11_robId,
  output wire [5:0]    io_contexts_11_euCtx_0,
  output wire [5:0]    io_contexts_11_euCtx_1,
  output wire [0:0]    io_contexts_12_staticWake,
  output wire [5:0]    io_contexts_12_physRd,
  output wire [5:0]    io_contexts_12_robId,
  output wire [5:0]    io_contexts_12_euCtx_0,
  output wire [5:0]    io_contexts_12_euCtx_1,
  output wire [0:0]    io_contexts_13_staticWake,
  output wire [5:0]    io_contexts_13_physRd,
  output wire [5:0]    io_contexts_13_robId,
  output wire [5:0]    io_contexts_13_euCtx_0,
  output wire [5:0]    io_contexts_13_euCtx_1,
  output wire [0:0]    io_contexts_14_staticWake,
  output wire [5:0]    io_contexts_14_physRd,
  output wire [5:0]    io_contexts_14_robId,
  output wire [5:0]    io_contexts_14_euCtx_0,
  output wire [5:0]    io_contexts_14_euCtx_1,
  output wire [0:0]    io_contexts_15_staticWake,
  output wire [5:0]    io_contexts_15_physRd,
  output wire [5:0]    io_contexts_15_robId,
  output wire [5:0]    io_contexts_15_euCtx_0,
  output wire [5:0]    io_contexts_15_euCtx_1,
  output wire [0:0]    io_contexts_16_staticWake,
  output wire [5:0]    io_contexts_16_physRd,
  output wire [5:0]    io_contexts_16_robId,
  output wire [5:0]    io_contexts_16_euCtx_0,
  output wire [5:0]    io_contexts_16_euCtx_1,
  output wire [0:0]    io_contexts_17_staticWake,
  output wire [5:0]    io_contexts_17_physRd,
  output wire [5:0]    io_contexts_17_robId,
  output wire [5:0]    io_contexts_17_euCtx_0,
  output wire [5:0]    io_contexts_17_euCtx_1,
  output wire [0:0]    io_contexts_18_staticWake,
  output wire [5:0]    io_contexts_18_physRd,
  output wire [5:0]    io_contexts_18_robId,
  output wire [5:0]    io_contexts_18_euCtx_0,
  output wire [5:0]    io_contexts_18_euCtx_1,
  output wire [0:0]    io_contexts_19_staticWake,
  output wire [5:0]    io_contexts_19_physRd,
  output wire [5:0]    io_contexts_19_robId,
  output wire [5:0]    io_contexts_19_euCtx_0,
  output wire [5:0]    io_contexts_19_euCtx_1,
  output wire [0:0]    io_contexts_20_staticWake,
  output wire [5:0]    io_contexts_20_physRd,
  output wire [5:0]    io_contexts_20_robId,
  output wire [5:0]    io_contexts_20_euCtx_0,
  output wire [5:0]    io_contexts_20_euCtx_1,
  output wire [0:0]    io_contexts_21_staticWake,
  output wire [5:0]    io_contexts_21_physRd,
  output wire [5:0]    io_contexts_21_robId,
  output wire [5:0]    io_contexts_21_euCtx_0,
  output wire [5:0]    io_contexts_21_euCtx_1,
  output wire [0:0]    io_contexts_22_staticWake,
  output wire [5:0]    io_contexts_22_physRd,
  output wire [5:0]    io_contexts_22_robId,
  output wire [5:0]    io_contexts_22_euCtx_0,
  output wire [5:0]    io_contexts_22_euCtx_1,
  output wire [0:0]    io_contexts_23_staticWake,
  output wire [5:0]    io_contexts_23_physRd,
  output wire [5:0]    io_contexts_23_robId,
  output wire [5:0]    io_contexts_23_euCtx_0,
  output wire [5:0]    io_contexts_23_euCtx_1,
  output wire [0:0]    io_contexts_24_staticWake,
  output wire [5:0]    io_contexts_24_physRd,
  output wire [5:0]    io_contexts_24_robId,
  output wire [5:0]    io_contexts_24_euCtx_0,
  output wire [5:0]    io_contexts_24_euCtx_1,
  output wire [0:0]    io_contexts_25_staticWake,
  output wire [5:0]    io_contexts_25_physRd,
  output wire [5:0]    io_contexts_25_robId,
  output wire [5:0]    io_contexts_25_euCtx_0,
  output wire [5:0]    io_contexts_25_euCtx_1,
  output wire [0:0]    io_contexts_26_staticWake,
  output wire [5:0]    io_contexts_26_physRd,
  output wire [5:0]    io_contexts_26_robId,
  output wire [5:0]    io_contexts_26_euCtx_0,
  output wire [5:0]    io_contexts_26_euCtx_1,
  output wire [0:0]    io_contexts_27_staticWake,
  output wire [5:0]    io_contexts_27_physRd,
  output wire [5:0]    io_contexts_27_robId,
  output wire [5:0]    io_contexts_27_euCtx_0,
  output wire [5:0]    io_contexts_27_euCtx_1,
  output wire [0:0]    io_contexts_28_staticWake,
  output wire [5:0]    io_contexts_28_physRd,
  output wire [5:0]    io_contexts_28_robId,
  output wire [5:0]    io_contexts_28_euCtx_0,
  output wire [5:0]    io_contexts_28_euCtx_1,
  output wire [0:0]    io_contexts_29_staticWake,
  output wire [5:0]    io_contexts_29_physRd,
  output wire [5:0]    io_contexts_29_robId,
  output wire [5:0]    io_contexts_29_euCtx_0,
  output wire [5:0]    io_contexts_29_euCtx_1,
  output wire [0:0]    io_contexts_30_staticWake,
  output wire [5:0]    io_contexts_30_physRd,
  output wire [5:0]    io_contexts_30_robId,
  output wire [5:0]    io_contexts_30_euCtx_0,
  output wire [5:0]    io_contexts_30_euCtx_1,
  output wire [0:0]    io_contexts_31_staticWake,
  output wire [5:0]    io_contexts_31_physRd,
  output wire [5:0]    io_contexts_31_robId,
  output wire [5:0]    io_contexts_31_euCtx_0,
  output wire [5:0]    io_contexts_31_euCtx_1,
  output reg  [31:0]   io_usage,
  input  wire          clk,
  input  wire          reset
);

  wire       [31:0]   _zz_event_moved;
  wire                _zz_selector_0_slotsValid;
  wire                _zz_selector_0_slotsValid_1;
  wire       [0:0]    _zz_selector_0_slotsValid_2;
  wire       [8:0]    _zz_selector_0_slotsValid_3;
  wire                _zz_selector_0_slotsValid_4;
  wire                _zz_selector_0_slotsValid_5;
  wire       [0:0]    _zz_selector_0_slotsValid_6;
  wire       [2:0]    _zz_selector_0_slotsValid_7;
  wire                _zz_selector_1_slotsValid;
  wire                _zz_selector_1_slotsValid_1;
  wire       [0:0]    _zz_selector_1_slotsValid_2;
  wire       [8:0]    _zz_selector_1_slotsValid_3;
  wire                _zz_selector_1_slotsValid_4;
  wire                _zz_selector_1_slotsValid_5;
  wire       [0:0]    _zz_selector_1_slotsValid_6;
  wire       [2:0]    _zz_selector_1_slotsValid_7;
  wire                _zz_selector_2_slotsValid;
  wire                _zz_selector_2_slotsValid_1;
  wire       [0:0]    _zz_selector_2_slotsValid_2;
  wire       [24:0]   _zz_selector_2_slotsValid_3;
  wire                _zz_selector_2_slotsValid_4;
  wire                _zz_selector_2_slotsValid_5;
  wire       [0:0]    _zz_selector_2_slotsValid_6;
  wire       [18:0]   _zz_selector_2_slotsValid_7;
  wire                _zz_selector_2_slotsValid_8;
  wire                _zz_selector_2_slotsValid_9;
  wire       [0:0]    _zz_selector_2_slotsValid_10;
  wire       [12:0]   _zz_selector_2_slotsValid_11;
  wire                _zz_selector_2_slotsValid_12;
  wire                _zz_selector_2_slotsValid_13;
  wire       [0:0]    _zz_selector_2_slotsValid_14;
  wire       [6:0]    _zz_selector_2_slotsValid_15;
  wire                _zz_selector_2_slotsValid_16;
  wire                _zz_selector_2_slotsValid_17;
  wire       [0:0]    _zz_selector_2_slotsValid_18;
  wire       [0:0]    _zz_selector_2_slotsValid_19;
  reg                 running;
  wire                clear;
  wire                lines_0_ways_0_fire;
  reg        [1:0]    lines_0_ways_0_sel;
  reg        [1:0]    lines_0_ways_0_selComb;
  reg        [0:0]    lines_0_ways_0_triggers;
  wire                lines_0_ways_0_ready;
  reg        [0:0]    lines_0_ways_0_context_staticWake;
  reg        [5:0]    lines_0_ways_0_context_physRd;
  reg        [5:0]    lines_0_ways_0_context_robId;
  reg        [5:0]    lines_0_ways_0_context_euCtx_0;
  reg        [5:0]    lines_0_ways_0_context_euCtx_1;
  wire                lines_0_ways_1_fire;
  reg        [1:0]    lines_0_ways_1_sel;
  reg        [1:0]    lines_0_ways_1_selComb;
  reg        [1:0]    lines_0_ways_1_triggers;
  wire                lines_0_ways_1_ready;
  reg        [0:0]    lines_0_ways_1_context_staticWake;
  reg        [5:0]    lines_0_ways_1_context_physRd;
  reg        [5:0]    lines_0_ways_1_context_robId;
  reg        [5:0]    lines_0_ways_1_context_euCtx_0;
  reg        [5:0]    lines_0_ways_1_context_euCtx_1;
  wire                lines_1_ways_0_fire;
  reg        [1:0]    lines_1_ways_0_sel;
  reg        [1:0]    lines_1_ways_0_selComb;
  reg        [2:0]    lines_1_ways_0_triggers;
  wire                lines_1_ways_0_ready;
  reg        [0:0]    lines_1_ways_0_context_staticWake;
  reg        [5:0]    lines_1_ways_0_context_physRd;
  reg        [5:0]    lines_1_ways_0_context_robId;
  reg        [5:0]    lines_1_ways_0_context_euCtx_0;
  reg        [5:0]    lines_1_ways_0_context_euCtx_1;
  wire                lines_1_ways_1_fire;
  reg        [1:0]    lines_1_ways_1_sel;
  reg        [1:0]    lines_1_ways_1_selComb;
  reg        [3:0]    lines_1_ways_1_triggers;
  wire                lines_1_ways_1_ready;
  reg        [0:0]    lines_1_ways_1_context_staticWake;
  reg        [5:0]    lines_1_ways_1_context_physRd;
  reg        [5:0]    lines_1_ways_1_context_robId;
  reg        [5:0]    lines_1_ways_1_context_euCtx_0;
  reg        [5:0]    lines_1_ways_1_context_euCtx_1;
  wire                lines_2_ways_0_fire;
  reg        [1:0]    lines_2_ways_0_sel;
  reg        [1:0]    lines_2_ways_0_selComb;
  reg        [4:0]    lines_2_ways_0_triggers;
  wire                lines_2_ways_0_ready;
  reg        [0:0]    lines_2_ways_0_context_staticWake;
  reg        [5:0]    lines_2_ways_0_context_physRd;
  reg        [5:0]    lines_2_ways_0_context_robId;
  reg        [5:0]    lines_2_ways_0_context_euCtx_0;
  reg        [5:0]    lines_2_ways_0_context_euCtx_1;
  wire                lines_2_ways_1_fire;
  reg        [1:0]    lines_2_ways_1_sel;
  reg        [1:0]    lines_2_ways_1_selComb;
  reg        [5:0]    lines_2_ways_1_triggers;
  wire                lines_2_ways_1_ready;
  reg        [0:0]    lines_2_ways_1_context_staticWake;
  reg        [5:0]    lines_2_ways_1_context_physRd;
  reg        [5:0]    lines_2_ways_1_context_robId;
  reg        [5:0]    lines_2_ways_1_context_euCtx_0;
  reg        [5:0]    lines_2_ways_1_context_euCtx_1;
  wire                lines_3_ways_0_fire;
  reg        [1:0]    lines_3_ways_0_sel;
  reg        [1:0]    lines_3_ways_0_selComb;
  reg        [6:0]    lines_3_ways_0_triggers;
  wire                lines_3_ways_0_ready;
  reg        [0:0]    lines_3_ways_0_context_staticWake;
  reg        [5:0]    lines_3_ways_0_context_physRd;
  reg        [5:0]    lines_3_ways_0_context_robId;
  reg        [5:0]    lines_3_ways_0_context_euCtx_0;
  reg        [5:0]    lines_3_ways_0_context_euCtx_1;
  wire                lines_3_ways_1_fire;
  reg        [1:0]    lines_3_ways_1_sel;
  reg        [1:0]    lines_3_ways_1_selComb;
  reg        [7:0]    lines_3_ways_1_triggers;
  wire                lines_3_ways_1_ready;
  reg        [0:0]    lines_3_ways_1_context_staticWake;
  reg        [5:0]    lines_3_ways_1_context_physRd;
  reg        [5:0]    lines_3_ways_1_context_robId;
  reg        [5:0]    lines_3_ways_1_context_euCtx_0;
  reg        [5:0]    lines_3_ways_1_context_euCtx_1;
  wire                lines_4_ways_0_fire;
  reg        [1:0]    lines_4_ways_0_sel;
  reg        [1:0]    lines_4_ways_0_selComb;
  reg        [8:0]    lines_4_ways_0_triggers;
  wire                lines_4_ways_0_ready;
  reg        [0:0]    lines_4_ways_0_context_staticWake;
  reg        [5:0]    lines_4_ways_0_context_physRd;
  reg        [5:0]    lines_4_ways_0_context_robId;
  reg        [5:0]    lines_4_ways_0_context_euCtx_0;
  reg        [5:0]    lines_4_ways_0_context_euCtx_1;
  wire                lines_4_ways_1_fire;
  reg        [1:0]    lines_4_ways_1_sel;
  reg        [1:0]    lines_4_ways_1_selComb;
  reg        [9:0]    lines_4_ways_1_triggers;
  wire                lines_4_ways_1_ready;
  reg        [0:0]    lines_4_ways_1_context_staticWake;
  reg        [5:0]    lines_4_ways_1_context_physRd;
  reg        [5:0]    lines_4_ways_1_context_robId;
  reg        [5:0]    lines_4_ways_1_context_euCtx_0;
  reg        [5:0]    lines_4_ways_1_context_euCtx_1;
  wire                lines_5_ways_0_fire;
  reg        [1:0]    lines_5_ways_0_sel;
  reg        [1:0]    lines_5_ways_0_selComb;
  reg        [10:0]   lines_5_ways_0_triggers;
  wire                lines_5_ways_0_ready;
  reg        [0:0]    lines_5_ways_0_context_staticWake;
  reg        [5:0]    lines_5_ways_0_context_physRd;
  reg        [5:0]    lines_5_ways_0_context_robId;
  reg        [5:0]    lines_5_ways_0_context_euCtx_0;
  reg        [5:0]    lines_5_ways_0_context_euCtx_1;
  wire                lines_5_ways_1_fire;
  reg        [1:0]    lines_5_ways_1_sel;
  reg        [1:0]    lines_5_ways_1_selComb;
  reg        [11:0]   lines_5_ways_1_triggers;
  wire                lines_5_ways_1_ready;
  reg        [0:0]    lines_5_ways_1_context_staticWake;
  reg        [5:0]    lines_5_ways_1_context_physRd;
  reg        [5:0]    lines_5_ways_1_context_robId;
  reg        [5:0]    lines_5_ways_1_context_euCtx_0;
  reg        [5:0]    lines_5_ways_1_context_euCtx_1;
  wire                lines_6_ways_0_fire;
  reg        [1:0]    lines_6_ways_0_sel;
  reg        [1:0]    lines_6_ways_0_selComb;
  reg        [12:0]   lines_6_ways_0_triggers;
  wire                lines_6_ways_0_ready;
  reg        [0:0]    lines_6_ways_0_context_staticWake;
  reg        [5:0]    lines_6_ways_0_context_physRd;
  reg        [5:0]    lines_6_ways_0_context_robId;
  reg        [5:0]    lines_6_ways_0_context_euCtx_0;
  reg        [5:0]    lines_6_ways_0_context_euCtx_1;
  wire                lines_6_ways_1_fire;
  reg        [1:0]    lines_6_ways_1_sel;
  reg        [1:0]    lines_6_ways_1_selComb;
  reg        [13:0]   lines_6_ways_1_triggers;
  wire                lines_6_ways_1_ready;
  reg        [0:0]    lines_6_ways_1_context_staticWake;
  reg        [5:0]    lines_6_ways_1_context_physRd;
  reg        [5:0]    lines_6_ways_1_context_robId;
  reg        [5:0]    lines_6_ways_1_context_euCtx_0;
  reg        [5:0]    lines_6_ways_1_context_euCtx_1;
  wire                lines_7_ways_0_fire;
  reg        [1:0]    lines_7_ways_0_sel;
  reg        [1:0]    lines_7_ways_0_selComb;
  reg        [14:0]   lines_7_ways_0_triggers;
  wire                lines_7_ways_0_ready;
  reg        [0:0]    lines_7_ways_0_context_staticWake;
  reg        [5:0]    lines_7_ways_0_context_physRd;
  reg        [5:0]    lines_7_ways_0_context_robId;
  reg        [5:0]    lines_7_ways_0_context_euCtx_0;
  reg        [5:0]    lines_7_ways_0_context_euCtx_1;
  wire                lines_7_ways_1_fire;
  reg        [1:0]    lines_7_ways_1_sel;
  reg        [1:0]    lines_7_ways_1_selComb;
  reg        [15:0]   lines_7_ways_1_triggers;
  wire                lines_7_ways_1_ready;
  reg        [0:0]    lines_7_ways_1_context_staticWake;
  reg        [5:0]    lines_7_ways_1_context_physRd;
  reg        [5:0]    lines_7_ways_1_context_robId;
  reg        [5:0]    lines_7_ways_1_context_euCtx_0;
  reg        [5:0]    lines_7_ways_1_context_euCtx_1;
  wire                lines_8_ways_0_fire;
  reg        [1:0]    lines_8_ways_0_sel;
  reg        [1:0]    lines_8_ways_0_selComb;
  reg        [16:0]   lines_8_ways_0_triggers;
  wire                lines_8_ways_0_ready;
  reg        [0:0]    lines_8_ways_0_context_staticWake;
  reg        [5:0]    lines_8_ways_0_context_physRd;
  reg        [5:0]    lines_8_ways_0_context_robId;
  reg        [5:0]    lines_8_ways_0_context_euCtx_0;
  reg        [5:0]    lines_8_ways_0_context_euCtx_1;
  wire                lines_8_ways_1_fire;
  reg        [1:0]    lines_8_ways_1_sel;
  reg        [1:0]    lines_8_ways_1_selComb;
  reg        [17:0]   lines_8_ways_1_triggers;
  wire                lines_8_ways_1_ready;
  reg        [0:0]    lines_8_ways_1_context_staticWake;
  reg        [5:0]    lines_8_ways_1_context_physRd;
  reg        [5:0]    lines_8_ways_1_context_robId;
  reg        [5:0]    lines_8_ways_1_context_euCtx_0;
  reg        [5:0]    lines_8_ways_1_context_euCtx_1;
  wire                lines_9_ways_0_fire;
  reg        [1:0]    lines_9_ways_0_sel;
  reg        [1:0]    lines_9_ways_0_selComb;
  reg        [18:0]   lines_9_ways_0_triggers;
  wire                lines_9_ways_0_ready;
  reg        [0:0]    lines_9_ways_0_context_staticWake;
  reg        [5:0]    lines_9_ways_0_context_physRd;
  reg        [5:0]    lines_9_ways_0_context_robId;
  reg        [5:0]    lines_9_ways_0_context_euCtx_0;
  reg        [5:0]    lines_9_ways_0_context_euCtx_1;
  wire                lines_9_ways_1_fire;
  reg        [1:0]    lines_9_ways_1_sel;
  reg        [1:0]    lines_9_ways_1_selComb;
  reg        [19:0]   lines_9_ways_1_triggers;
  wire                lines_9_ways_1_ready;
  reg        [0:0]    lines_9_ways_1_context_staticWake;
  reg        [5:0]    lines_9_ways_1_context_physRd;
  reg        [5:0]    lines_9_ways_1_context_robId;
  reg        [5:0]    lines_9_ways_1_context_euCtx_0;
  reg        [5:0]    lines_9_ways_1_context_euCtx_1;
  wire                lines_10_ways_0_fire;
  reg        [1:0]    lines_10_ways_0_sel;
  reg        [1:0]    lines_10_ways_0_selComb;
  reg        [20:0]   lines_10_ways_0_triggers;
  wire                lines_10_ways_0_ready;
  reg        [0:0]    lines_10_ways_0_context_staticWake;
  reg        [5:0]    lines_10_ways_0_context_physRd;
  reg        [5:0]    lines_10_ways_0_context_robId;
  reg        [5:0]    lines_10_ways_0_context_euCtx_0;
  reg        [5:0]    lines_10_ways_0_context_euCtx_1;
  wire                lines_10_ways_1_fire;
  reg        [1:0]    lines_10_ways_1_sel;
  reg        [1:0]    lines_10_ways_1_selComb;
  reg        [21:0]   lines_10_ways_1_triggers;
  wire                lines_10_ways_1_ready;
  reg        [0:0]    lines_10_ways_1_context_staticWake;
  reg        [5:0]    lines_10_ways_1_context_physRd;
  reg        [5:0]    lines_10_ways_1_context_robId;
  reg        [5:0]    lines_10_ways_1_context_euCtx_0;
  reg        [5:0]    lines_10_ways_1_context_euCtx_1;
  wire                lines_11_ways_0_fire;
  reg        [1:0]    lines_11_ways_0_sel;
  reg        [1:0]    lines_11_ways_0_selComb;
  reg        [22:0]   lines_11_ways_0_triggers;
  wire                lines_11_ways_0_ready;
  reg        [0:0]    lines_11_ways_0_context_staticWake;
  reg        [5:0]    lines_11_ways_0_context_physRd;
  reg        [5:0]    lines_11_ways_0_context_robId;
  reg        [5:0]    lines_11_ways_0_context_euCtx_0;
  reg        [5:0]    lines_11_ways_0_context_euCtx_1;
  wire                lines_11_ways_1_fire;
  reg        [1:0]    lines_11_ways_1_sel;
  reg        [1:0]    lines_11_ways_1_selComb;
  reg        [23:0]   lines_11_ways_1_triggers;
  wire                lines_11_ways_1_ready;
  reg        [0:0]    lines_11_ways_1_context_staticWake;
  reg        [5:0]    lines_11_ways_1_context_physRd;
  reg        [5:0]    lines_11_ways_1_context_robId;
  reg        [5:0]    lines_11_ways_1_context_euCtx_0;
  reg        [5:0]    lines_11_ways_1_context_euCtx_1;
  wire                lines_12_ways_0_fire;
  reg        [1:0]    lines_12_ways_0_sel;
  reg        [1:0]    lines_12_ways_0_selComb;
  reg        [24:0]   lines_12_ways_0_triggers;
  wire                lines_12_ways_0_ready;
  reg        [0:0]    lines_12_ways_0_context_staticWake;
  reg        [5:0]    lines_12_ways_0_context_physRd;
  reg        [5:0]    lines_12_ways_0_context_robId;
  reg        [5:0]    lines_12_ways_0_context_euCtx_0;
  reg        [5:0]    lines_12_ways_0_context_euCtx_1;
  wire                lines_12_ways_1_fire;
  reg        [1:0]    lines_12_ways_1_sel;
  reg        [1:0]    lines_12_ways_1_selComb;
  reg        [25:0]   lines_12_ways_1_triggers;
  wire                lines_12_ways_1_ready;
  reg        [0:0]    lines_12_ways_1_context_staticWake;
  reg        [5:0]    lines_12_ways_1_context_physRd;
  reg        [5:0]    lines_12_ways_1_context_robId;
  reg        [5:0]    lines_12_ways_1_context_euCtx_0;
  reg        [5:0]    lines_12_ways_1_context_euCtx_1;
  wire                lines_13_ways_0_fire;
  reg        [1:0]    lines_13_ways_0_sel;
  reg        [1:0]    lines_13_ways_0_selComb;
  reg        [26:0]   lines_13_ways_0_triggers;
  wire                lines_13_ways_0_ready;
  reg        [0:0]    lines_13_ways_0_context_staticWake;
  reg        [5:0]    lines_13_ways_0_context_physRd;
  reg        [5:0]    lines_13_ways_0_context_robId;
  reg        [5:0]    lines_13_ways_0_context_euCtx_0;
  reg        [5:0]    lines_13_ways_0_context_euCtx_1;
  wire                lines_13_ways_1_fire;
  reg        [1:0]    lines_13_ways_1_sel;
  reg        [1:0]    lines_13_ways_1_selComb;
  reg        [27:0]   lines_13_ways_1_triggers;
  wire                lines_13_ways_1_ready;
  reg        [0:0]    lines_13_ways_1_context_staticWake;
  reg        [5:0]    lines_13_ways_1_context_physRd;
  reg        [5:0]    lines_13_ways_1_context_robId;
  reg        [5:0]    lines_13_ways_1_context_euCtx_0;
  reg        [5:0]    lines_13_ways_1_context_euCtx_1;
  wire                lines_14_ways_0_fire;
  reg        [1:0]    lines_14_ways_0_sel;
  reg        [1:0]    lines_14_ways_0_selComb;
  reg        [28:0]   lines_14_ways_0_triggers;
  wire                lines_14_ways_0_ready;
  reg        [0:0]    lines_14_ways_0_context_staticWake;
  reg        [5:0]    lines_14_ways_0_context_physRd;
  reg        [5:0]    lines_14_ways_0_context_robId;
  reg        [5:0]    lines_14_ways_0_context_euCtx_0;
  reg        [5:0]    lines_14_ways_0_context_euCtx_1;
  wire                lines_14_ways_1_fire;
  reg        [1:0]    lines_14_ways_1_sel;
  reg        [1:0]    lines_14_ways_1_selComb;
  reg        [29:0]   lines_14_ways_1_triggers;
  wire                lines_14_ways_1_ready;
  reg        [0:0]    lines_14_ways_1_context_staticWake;
  reg        [5:0]    lines_14_ways_1_context_physRd;
  reg        [5:0]    lines_14_ways_1_context_robId;
  reg        [5:0]    lines_14_ways_1_context_euCtx_0;
  reg        [5:0]    lines_14_ways_1_context_euCtx_1;
  wire                lines_15_ways_0_fire;
  reg        [1:0]    lines_15_ways_0_sel;
  reg        [1:0]    lines_15_ways_0_selComb;
  reg        [30:0]   lines_15_ways_0_triggers;
  wire                lines_15_ways_0_ready;
  reg        [0:0]    lines_15_ways_0_context_staticWake;
  reg        [5:0]    lines_15_ways_0_context_physRd;
  reg        [5:0]    lines_15_ways_0_context_robId;
  reg        [5:0]    lines_15_ways_0_context_euCtx_0;
  reg        [5:0]    lines_15_ways_0_context_euCtx_1;
  wire                lines_15_ways_1_fire;
  reg        [1:0]    lines_15_ways_1_sel;
  reg        [1:0]    lines_15_ways_1_selComb;
  reg        [31:0]   lines_15_ways_1_triggers;
  wire                lines_15_ways_1_ready;
  reg        [0:0]    lines_15_ways_1_context_staticWake;
  reg        [5:0]    lines_15_ways_1_context_physRd;
  reg        [5:0]    lines_15_ways_1_context_robId;
  reg        [5:0]    lines_15_ways_1_context_euCtx_0;
  reg        [5:0]    lines_15_ways_1_context_euCtx_1;
  wire                compaction_moveIt;
  wire       [31:0]   event_moved;
  wire       [31:0]   event_value;
  wire                when_IssueQueue_l109;
  wire                when_IssueQueue_l109_1;
  wire                when_IssueQueue_l109_2;
  wire                when_IssueQueue_l109_3;
  wire                when_IssueQueue_l109_4;
  wire                when_IssueQueue_l109_5;
  wire                when_IssueQueue_l109_6;
  wire                when_IssueQueue_l109_7;
  wire                when_IssueQueue_l109_8;
  wire                when_IssueQueue_l109_9;
  wire                when_IssueQueue_l109_10;
  wire                when_IssueQueue_l109_11;
  wire                when_IssueQueue_l109_12;
  wire                when_IssueQueue_l109_13;
  wire                when_IssueQueue_l109_14;
  wire                when_IssueQueue_l109_15;
  wire                when_IssueQueue_l109_16;
  wire                when_IssueQueue_l109_17;
  wire                when_IssueQueue_l109_18;
  wire                when_IssueQueue_l109_19;
  wire                when_IssueQueue_l109_20;
  wire                when_IssueQueue_l109_21;
  wire                when_IssueQueue_l109_22;
  wire                when_IssueQueue_l109_23;
  wire                when_IssueQueue_l109_24;
  wire                when_IssueQueue_l109_25;
  wire                when_IssueQueue_l109_26;
  wire                when_IssueQueue_l109_27;
  wire                when_IssueQueue_l109_28;
  wire                when_IssueQueue_l109_29;
  wire                when_IssueQueue_l109_30;
  wire                when_IssueQueue_l109_31;
  wire       [15:0]   selector_0_slotsValid;
  wire       [15:0]   _zz_selector_0_slotsValid_bools_0;
  wire                selector_0_slotsValid_bools_0;
  wire                selector_0_slotsValid_bools_1;
  wire                selector_0_slotsValid_bools_2;
  wire                selector_0_slotsValid_bools_3;
  wire                selector_0_slotsValid_bools_4;
  wire                selector_0_slotsValid_bools_5;
  wire                selector_0_slotsValid_bools_6;
  wire                selector_0_slotsValid_bools_7;
  wire                selector_0_slotsValid_bools_8;
  wire                selector_0_slotsValid_bools_9;
  wire                selector_0_slotsValid_bools_10;
  wire                selector_0_slotsValid_bools_11;
  wire                selector_0_slotsValid_bools_12;
  wire                selector_0_slotsValid_bools_13;
  wire                selector_0_slotsValid_bools_14;
  wire                selector_0_slotsValid_bools_15;
  reg        [15:0]   _zz_selector_0_selOh;
  wire                selector_0_slotsValid_range_0_to_1;
  wire                selector_0_slotsValid_range_0_to_2;
  wire                selector_0_slotsValid_range_0_to_3;
  wire                selector_0_slotsValid_range_0_to_4;
  wire                selector_0_slotsValid_range_0_to_5;
  wire                selector_0_slotsValid_range_6_to_7;
  wire                selector_0_slotsValid_range_6_to_8;
  wire                selector_0_slotsValid_range_6_to_9;
  wire                selector_0_slotsValid_range_6_to_10;
  wire                selector_0_slotsValid_range_6_to_11;
  wire                selector_0_slotsValid_range_0_to_11;
  wire                selector_0_slotsValid_range_12_to_13;
  wire                selector_0_slotsValid_range_12_to_14;
  wire       [15:0]   selector_0_selOh;
  wire       [15:0]   selector_1_slotsValid;
  wire       [15:0]   _zz_selector_1_slotsValid_bools_0;
  wire                selector_1_slotsValid_bools_0;
  wire                selector_1_slotsValid_bools_1;
  wire                selector_1_slotsValid_bools_2;
  wire                selector_1_slotsValid_bools_3;
  wire                selector_1_slotsValid_bools_4;
  wire                selector_1_slotsValid_bools_5;
  wire                selector_1_slotsValid_bools_6;
  wire                selector_1_slotsValid_bools_7;
  wire                selector_1_slotsValid_bools_8;
  wire                selector_1_slotsValid_bools_9;
  wire                selector_1_slotsValid_bools_10;
  wire                selector_1_slotsValid_bools_11;
  wire                selector_1_slotsValid_bools_12;
  wire                selector_1_slotsValid_bools_13;
  wire                selector_1_slotsValid_bools_14;
  wire                selector_1_slotsValid_bools_15;
  reg        [15:0]   _zz_selector_1_selOh;
  wire                selector_1_slotsValid_range_0_to_1;
  wire                selector_1_slotsValid_range_0_to_2;
  wire                selector_1_slotsValid_range_0_to_3;
  wire                selector_1_slotsValid_range_0_to_4;
  wire                selector_1_slotsValid_range_0_to_5;
  wire                selector_1_slotsValid_range_6_to_7;
  wire                selector_1_slotsValid_range_6_to_8;
  wire                selector_1_slotsValid_range_6_to_9;
  wire                selector_1_slotsValid_range_6_to_10;
  wire                selector_1_slotsValid_range_6_to_11;
  wire                selector_1_slotsValid_range_0_to_11;
  wire                selector_1_slotsValid_range_12_to_13;
  wire                selector_1_slotsValid_range_12_to_14;
  wire       [15:0]   selector_1_selOh;
  wire       [31:0]   selector_2_slotsValid;
  wire       [31:0]   _zz_selector_2_slotsValid_bools_0;
  wire                selector_2_slotsValid_bools_0;
  wire                selector_2_slotsValid_bools_1;
  wire                selector_2_slotsValid_bools_2;
  wire                selector_2_slotsValid_bools_3;
  wire                selector_2_slotsValid_bools_4;
  wire                selector_2_slotsValid_bools_5;
  wire                selector_2_slotsValid_bools_6;
  wire                selector_2_slotsValid_bools_7;
  wire                selector_2_slotsValid_bools_8;
  wire                selector_2_slotsValid_bools_9;
  wire                selector_2_slotsValid_bools_10;
  wire                selector_2_slotsValid_bools_11;
  wire                selector_2_slotsValid_bools_12;
  wire                selector_2_slotsValid_bools_13;
  wire                selector_2_slotsValid_bools_14;
  wire                selector_2_slotsValid_bools_15;
  wire                selector_2_slotsValid_bools_16;
  wire                selector_2_slotsValid_bools_17;
  wire                selector_2_slotsValid_bools_18;
  wire                selector_2_slotsValid_bools_19;
  wire                selector_2_slotsValid_bools_20;
  wire                selector_2_slotsValid_bools_21;
  wire                selector_2_slotsValid_bools_22;
  wire                selector_2_slotsValid_bools_23;
  wire                selector_2_slotsValid_bools_24;
  wire                selector_2_slotsValid_bools_25;
  wire                selector_2_slotsValid_bools_26;
  wire                selector_2_slotsValid_bools_27;
  wire                selector_2_slotsValid_bools_28;
  wire                selector_2_slotsValid_bools_29;
  wire                selector_2_slotsValid_bools_30;
  wire                selector_2_slotsValid_bools_31;
  reg        [31:0]   _zz_selector_2_selOh;
  wire                selector_2_slotsValid_range_0_to_1;
  wire                selector_2_slotsValid_range_0_to_2;
  wire                selector_2_slotsValid_range_0_to_3;
  wire                selector_2_slotsValid_range_0_to_4;
  wire                selector_2_slotsValid_range_0_to_5;
  wire                selector_2_slotsValid_range_6_to_7;
  wire                selector_2_slotsValid_range_6_to_8;
  wire                selector_2_slotsValid_range_6_to_9;
  wire                selector_2_slotsValid_range_6_to_10;
  wire                selector_2_slotsValid_range_6_to_11;
  wire                selector_2_slotsValid_range_0_to_11;
  wire                selector_2_slotsValid_range_12_to_13;
  wire                selector_2_slotsValid_range_12_to_14;
  wire                selector_2_slotsValid_range_12_to_15;
  wire                selector_2_slotsValid_range_12_to_16;
  wire                selector_2_slotsValid_range_12_to_17;
  wire                selector_2_slotsValid_range_0_to_17;
  wire                selector_2_slotsValid_range_18_to_19;
  wire                selector_2_slotsValid_range_18_to_20;
  wire                selector_2_slotsValid_range_18_to_21;
  wire                selector_2_slotsValid_range_18_to_22;
  wire                selector_2_slotsValid_range_18_to_23;
  wire                selector_2_slotsValid_range_0_to_23;
  wire                selector_2_slotsValid_range_24_to_25;
  wire                selector_2_slotsValid_range_24_to_26;
  wire                selector_2_slotsValid_range_24_to_27;
  wire                selector_2_slotsValid_range_24_to_28;
  wire                selector_2_slotsValid_range_24_to_29;
  wire                selector_2_slotsValid_range_0_to_29;
  wire       [31:0]   selector_2_selOh;
  wire                line0Ready;
  wire                line1Ready;
  reg                 readyReg;

  assign _zz_event_moved = (io_events >>> 2);
  assign _zz_selector_0_slotsValid = lines_11_ways_0_sel[0];
  assign _zz_selector_0_slotsValid_1 = (lines_10_ways_0_ready && lines_10_ways_0_sel[0]);
  assign _zz_selector_0_slotsValid_2 = (lines_9_ways_0_ready && lines_9_ways_0_sel[0]);
  assign _zz_selector_0_slotsValid_3 = {(lines_8_ways_0_ready && lines_8_ways_0_sel[0]),{(lines_7_ways_0_ready && lines_7_ways_0_sel[0]),{(lines_6_ways_0_ready && lines_6_ways_0_sel[0]),{(lines_5_ways_0_ready && _zz_selector_0_slotsValid_4),{_zz_selector_0_slotsValid_5,{_zz_selector_0_slotsValid_6,_zz_selector_0_slotsValid_7}}}}}};
  assign _zz_selector_0_slotsValid_4 = lines_5_ways_0_sel[0];
  assign _zz_selector_0_slotsValid_5 = (lines_4_ways_0_ready && lines_4_ways_0_sel[0]);
  assign _zz_selector_0_slotsValid_6 = (lines_3_ways_0_ready && lines_3_ways_0_sel[0]);
  assign _zz_selector_0_slotsValid_7 = {(lines_2_ways_0_ready && lines_2_ways_0_sel[0]),{(lines_1_ways_0_ready && lines_1_ways_0_sel[0]),(lines_0_ways_0_ready && lines_0_ways_0_sel[0])}};
  assign _zz_selector_1_slotsValid = lines_11_ways_1_sel[0];
  assign _zz_selector_1_slotsValid_1 = (lines_10_ways_1_ready && lines_10_ways_1_sel[0]);
  assign _zz_selector_1_slotsValid_2 = (lines_9_ways_1_ready && lines_9_ways_1_sel[0]);
  assign _zz_selector_1_slotsValid_3 = {(lines_8_ways_1_ready && lines_8_ways_1_sel[0]),{(lines_7_ways_1_ready && lines_7_ways_1_sel[0]),{(lines_6_ways_1_ready && lines_6_ways_1_sel[0]),{(lines_5_ways_1_ready && _zz_selector_1_slotsValid_4),{_zz_selector_1_slotsValid_5,{_zz_selector_1_slotsValid_6,_zz_selector_1_slotsValid_7}}}}}};
  assign _zz_selector_1_slotsValid_4 = lines_5_ways_1_sel[0];
  assign _zz_selector_1_slotsValid_5 = (lines_4_ways_1_ready && lines_4_ways_1_sel[0]);
  assign _zz_selector_1_slotsValid_6 = (lines_3_ways_1_ready && lines_3_ways_1_sel[0]);
  assign _zz_selector_1_slotsValid_7 = {(lines_2_ways_1_ready && lines_2_ways_1_sel[0]),{(lines_1_ways_1_ready && lines_1_ways_1_sel[0]),(lines_0_ways_1_ready && lines_0_ways_1_sel[0])}};
  assign _zz_selector_2_slotsValid = lines_13_ways_1_sel[1];
  assign _zz_selector_2_slotsValid_1 = (lines_13_ways_0_ready && lines_13_ways_0_sel[1]);
  assign _zz_selector_2_slotsValid_2 = (lines_12_ways_1_ready && lines_12_ways_1_sel[1]);
  assign _zz_selector_2_slotsValid_3 = {(lines_12_ways_0_ready && lines_12_ways_0_sel[1]),{(lines_11_ways_1_ready && lines_11_ways_1_sel[1]),{(lines_11_ways_0_ready && lines_11_ways_0_sel[1]),{(lines_10_ways_1_ready && _zz_selector_2_slotsValid_4),{_zz_selector_2_slotsValid_5,{_zz_selector_2_slotsValid_6,_zz_selector_2_slotsValid_7}}}}}};
  assign _zz_selector_2_slotsValid_4 = lines_10_ways_1_sel[1];
  assign _zz_selector_2_slotsValid_5 = (lines_10_ways_0_ready && lines_10_ways_0_sel[1]);
  assign _zz_selector_2_slotsValid_6 = (lines_9_ways_1_ready && lines_9_ways_1_sel[1]);
  assign _zz_selector_2_slotsValid_7 = {(lines_9_ways_0_ready && lines_9_ways_0_sel[1]),{(lines_8_ways_1_ready && lines_8_ways_1_sel[1]),{(lines_8_ways_0_ready && lines_8_ways_0_sel[1]),{(lines_7_ways_1_ready && _zz_selector_2_slotsValid_8),{_zz_selector_2_slotsValid_9,{_zz_selector_2_slotsValid_10,_zz_selector_2_slotsValid_11}}}}}};
  assign _zz_selector_2_slotsValid_8 = lines_7_ways_1_sel[1];
  assign _zz_selector_2_slotsValid_9 = (lines_7_ways_0_ready && lines_7_ways_0_sel[1]);
  assign _zz_selector_2_slotsValid_10 = (lines_6_ways_1_ready && lines_6_ways_1_sel[1]);
  assign _zz_selector_2_slotsValid_11 = {(lines_6_ways_0_ready && lines_6_ways_0_sel[1]),{(lines_5_ways_1_ready && lines_5_ways_1_sel[1]),{(lines_5_ways_0_ready && lines_5_ways_0_sel[1]),{(lines_4_ways_1_ready && _zz_selector_2_slotsValid_12),{_zz_selector_2_slotsValid_13,{_zz_selector_2_slotsValid_14,_zz_selector_2_slotsValid_15}}}}}};
  assign _zz_selector_2_slotsValid_12 = lines_4_ways_1_sel[1];
  assign _zz_selector_2_slotsValid_13 = (lines_4_ways_0_ready && lines_4_ways_0_sel[1]);
  assign _zz_selector_2_slotsValid_14 = (lines_3_ways_1_ready && lines_3_ways_1_sel[1]);
  assign _zz_selector_2_slotsValid_15 = {(lines_3_ways_0_ready && lines_3_ways_0_sel[1]),{(lines_2_ways_1_ready && lines_2_ways_1_sel[1]),{(lines_2_ways_0_ready && lines_2_ways_0_sel[1]),{(lines_1_ways_1_ready && _zz_selector_2_slotsValid_16),{_zz_selector_2_slotsValid_17,{_zz_selector_2_slotsValid_18,_zz_selector_2_slotsValid_19}}}}}};
  assign _zz_selector_2_slotsValid_16 = lines_1_ways_1_sel[1];
  assign _zz_selector_2_slotsValid_17 = (lines_1_ways_0_ready && lines_1_ways_0_sel[1]);
  assign _zz_selector_2_slotsValid_18 = (lines_0_ways_1_ready && lines_0_ways_1_sel[1]);
  assign _zz_selector_2_slotsValid_19 = (lines_0_ways_0_ready && lines_0_ways_0_sel[1]);
  assign clear = (io_clear || (! running));
  always @(*) begin
    lines_0_ways_0_selComb = lines_0_ways_0_sel;
    if(lines_0_ways_0_fire) begin
      lines_0_ways_0_selComb = 2'b00;
    end
  end

  assign lines_0_ways_0_ready = 1'b1;
  assign io_contexts_0_staticWake = lines_0_ways_0_context_staticWake;
  assign io_contexts_0_physRd = lines_0_ways_0_context_physRd;
  assign io_contexts_0_robId = lines_0_ways_0_context_robId;
  assign io_contexts_0_euCtx_0 = lines_0_ways_0_context_euCtx_0;
  assign io_contexts_0_euCtx_1 = lines_0_ways_0_context_euCtx_1;
  always @(*) begin
    io_usage[0] = ((lines_0_ways_0_sel != 2'b00) || lines_0_ways_0_triggers[0]);
    io_usage[1] = ((lines_0_ways_1_sel != 2'b00) || lines_0_ways_1_triggers[1]);
    io_usage[2] = ((lines_1_ways_0_sel != 2'b00) || lines_1_ways_0_triggers[2]);
    io_usage[3] = ((lines_1_ways_1_sel != 2'b00) || lines_1_ways_1_triggers[3]);
    io_usage[4] = ((lines_2_ways_0_sel != 2'b00) || lines_2_ways_0_triggers[4]);
    io_usage[5] = ((lines_2_ways_1_sel != 2'b00) || lines_2_ways_1_triggers[5]);
    io_usage[6] = ((lines_3_ways_0_sel != 2'b00) || lines_3_ways_0_triggers[6]);
    io_usage[7] = ((lines_3_ways_1_sel != 2'b00) || lines_3_ways_1_triggers[7]);
    io_usage[8] = ((lines_4_ways_0_sel != 2'b00) || lines_4_ways_0_triggers[8]);
    io_usage[9] = ((lines_4_ways_1_sel != 2'b00) || lines_4_ways_1_triggers[9]);
    io_usage[10] = ((lines_5_ways_0_sel != 2'b00) || lines_5_ways_0_triggers[10]);
    io_usage[11] = ((lines_5_ways_1_sel != 2'b00) || lines_5_ways_1_triggers[11]);
    io_usage[12] = ((lines_6_ways_0_sel != 2'b00) || lines_6_ways_0_triggers[12]);
    io_usage[13] = ((lines_6_ways_1_sel != 2'b00) || lines_6_ways_1_triggers[13]);
    io_usage[14] = ((lines_7_ways_0_sel != 2'b00) || lines_7_ways_0_triggers[14]);
    io_usage[15] = ((lines_7_ways_1_sel != 2'b00) || lines_7_ways_1_triggers[15]);
    io_usage[16] = ((lines_8_ways_0_sel != 2'b00) || lines_8_ways_0_triggers[16]);
    io_usage[17] = ((lines_8_ways_1_sel != 2'b00) || lines_8_ways_1_triggers[17]);
    io_usage[18] = ((lines_9_ways_0_sel != 2'b00) || lines_9_ways_0_triggers[18]);
    io_usage[19] = ((lines_9_ways_1_sel != 2'b00) || lines_9_ways_1_triggers[19]);
    io_usage[20] = ((lines_10_ways_0_sel != 2'b00) || lines_10_ways_0_triggers[20]);
    io_usage[21] = ((lines_10_ways_1_sel != 2'b00) || lines_10_ways_1_triggers[21]);
    io_usage[22] = ((lines_11_ways_0_sel != 2'b00) || lines_11_ways_0_triggers[22]);
    io_usage[23] = ((lines_11_ways_1_sel != 2'b00) || lines_11_ways_1_triggers[23]);
    io_usage[24] = ((lines_12_ways_0_sel != 2'b00) || lines_12_ways_0_triggers[24]);
    io_usage[25] = ((lines_12_ways_1_sel != 2'b00) || lines_12_ways_1_triggers[25]);
    io_usage[26] = ((lines_13_ways_0_sel != 2'b00) || lines_13_ways_0_triggers[26]);
    io_usage[27] = ((lines_13_ways_1_sel != 2'b00) || lines_13_ways_1_triggers[27]);
    io_usage[28] = ((lines_14_ways_0_sel != 2'b00) || lines_14_ways_0_triggers[28]);
    io_usage[29] = ((lines_14_ways_1_sel != 2'b00) || lines_14_ways_1_triggers[29]);
    io_usage[30] = ((lines_15_ways_0_sel != 2'b00) || lines_15_ways_0_triggers[30]);
    io_usage[31] = ((lines_15_ways_1_sel != 2'b00) || lines_15_ways_1_triggers[31]);
  end

  always @(*) begin
    lines_0_ways_1_selComb = lines_0_ways_1_sel;
    if(lines_0_ways_1_fire) begin
      lines_0_ways_1_selComb = 2'b00;
    end
  end

  assign lines_0_ways_1_ready = (lines_0_ways_1_triggers[0 : 0] == 1'b0);
  assign io_contexts_1_staticWake = lines_0_ways_1_context_staticWake;
  assign io_contexts_1_physRd = lines_0_ways_1_context_physRd;
  assign io_contexts_1_robId = lines_0_ways_1_context_robId;
  assign io_contexts_1_euCtx_0 = lines_0_ways_1_context_euCtx_0;
  assign io_contexts_1_euCtx_1 = lines_0_ways_1_context_euCtx_1;
  always @(*) begin
    lines_1_ways_0_selComb = lines_1_ways_0_sel;
    if(lines_1_ways_0_fire) begin
      lines_1_ways_0_selComb = 2'b00;
    end
  end

  assign lines_1_ways_0_ready = (lines_1_ways_0_triggers[1 : 0] == 2'b00);
  assign io_contexts_2_staticWake = lines_1_ways_0_context_staticWake;
  assign io_contexts_2_physRd = lines_1_ways_0_context_physRd;
  assign io_contexts_2_robId = lines_1_ways_0_context_robId;
  assign io_contexts_2_euCtx_0 = lines_1_ways_0_context_euCtx_0;
  assign io_contexts_2_euCtx_1 = lines_1_ways_0_context_euCtx_1;
  always @(*) begin
    lines_1_ways_1_selComb = lines_1_ways_1_sel;
    if(lines_1_ways_1_fire) begin
      lines_1_ways_1_selComb = 2'b00;
    end
  end

  assign lines_1_ways_1_ready = (lines_1_ways_1_triggers[2 : 0] == 3'b000);
  assign io_contexts_3_staticWake = lines_1_ways_1_context_staticWake;
  assign io_contexts_3_physRd = lines_1_ways_1_context_physRd;
  assign io_contexts_3_robId = lines_1_ways_1_context_robId;
  assign io_contexts_3_euCtx_0 = lines_1_ways_1_context_euCtx_0;
  assign io_contexts_3_euCtx_1 = lines_1_ways_1_context_euCtx_1;
  always @(*) begin
    lines_2_ways_0_selComb = lines_2_ways_0_sel;
    if(lines_2_ways_0_fire) begin
      lines_2_ways_0_selComb = 2'b00;
    end
  end

  assign lines_2_ways_0_ready = (lines_2_ways_0_triggers[3 : 0] == 4'b0000);
  assign io_contexts_4_staticWake = lines_2_ways_0_context_staticWake;
  assign io_contexts_4_physRd = lines_2_ways_0_context_physRd;
  assign io_contexts_4_robId = lines_2_ways_0_context_robId;
  assign io_contexts_4_euCtx_0 = lines_2_ways_0_context_euCtx_0;
  assign io_contexts_4_euCtx_1 = lines_2_ways_0_context_euCtx_1;
  always @(*) begin
    lines_2_ways_1_selComb = lines_2_ways_1_sel;
    if(lines_2_ways_1_fire) begin
      lines_2_ways_1_selComb = 2'b00;
    end
  end

  assign lines_2_ways_1_ready = (lines_2_ways_1_triggers[4 : 0] == 5'h00);
  assign io_contexts_5_staticWake = lines_2_ways_1_context_staticWake;
  assign io_contexts_5_physRd = lines_2_ways_1_context_physRd;
  assign io_contexts_5_robId = lines_2_ways_1_context_robId;
  assign io_contexts_5_euCtx_0 = lines_2_ways_1_context_euCtx_0;
  assign io_contexts_5_euCtx_1 = lines_2_ways_1_context_euCtx_1;
  always @(*) begin
    lines_3_ways_0_selComb = lines_3_ways_0_sel;
    if(lines_3_ways_0_fire) begin
      lines_3_ways_0_selComb = 2'b00;
    end
  end

  assign lines_3_ways_0_ready = (lines_3_ways_0_triggers[5 : 0] == 6'h00);
  assign io_contexts_6_staticWake = lines_3_ways_0_context_staticWake;
  assign io_contexts_6_physRd = lines_3_ways_0_context_physRd;
  assign io_contexts_6_robId = lines_3_ways_0_context_robId;
  assign io_contexts_6_euCtx_0 = lines_3_ways_0_context_euCtx_0;
  assign io_contexts_6_euCtx_1 = lines_3_ways_0_context_euCtx_1;
  always @(*) begin
    lines_3_ways_1_selComb = lines_3_ways_1_sel;
    if(lines_3_ways_1_fire) begin
      lines_3_ways_1_selComb = 2'b00;
    end
  end

  assign lines_3_ways_1_ready = (lines_3_ways_1_triggers[6 : 0] == 7'h00);
  assign io_contexts_7_staticWake = lines_3_ways_1_context_staticWake;
  assign io_contexts_7_physRd = lines_3_ways_1_context_physRd;
  assign io_contexts_7_robId = lines_3_ways_1_context_robId;
  assign io_contexts_7_euCtx_0 = lines_3_ways_1_context_euCtx_0;
  assign io_contexts_7_euCtx_1 = lines_3_ways_1_context_euCtx_1;
  always @(*) begin
    lines_4_ways_0_selComb = lines_4_ways_0_sel;
    if(lines_4_ways_0_fire) begin
      lines_4_ways_0_selComb = 2'b00;
    end
  end

  assign lines_4_ways_0_ready = (lines_4_ways_0_triggers[7 : 0] == 8'h00);
  assign io_contexts_8_staticWake = lines_4_ways_0_context_staticWake;
  assign io_contexts_8_physRd = lines_4_ways_0_context_physRd;
  assign io_contexts_8_robId = lines_4_ways_0_context_robId;
  assign io_contexts_8_euCtx_0 = lines_4_ways_0_context_euCtx_0;
  assign io_contexts_8_euCtx_1 = lines_4_ways_0_context_euCtx_1;
  always @(*) begin
    lines_4_ways_1_selComb = lines_4_ways_1_sel;
    if(lines_4_ways_1_fire) begin
      lines_4_ways_1_selComb = 2'b00;
    end
  end

  assign lines_4_ways_1_ready = (lines_4_ways_1_triggers[8 : 0] == 9'h000);
  assign io_contexts_9_staticWake = lines_4_ways_1_context_staticWake;
  assign io_contexts_9_physRd = lines_4_ways_1_context_physRd;
  assign io_contexts_9_robId = lines_4_ways_1_context_robId;
  assign io_contexts_9_euCtx_0 = lines_4_ways_1_context_euCtx_0;
  assign io_contexts_9_euCtx_1 = lines_4_ways_1_context_euCtx_1;
  always @(*) begin
    lines_5_ways_0_selComb = lines_5_ways_0_sel;
    if(lines_5_ways_0_fire) begin
      lines_5_ways_0_selComb = 2'b00;
    end
  end

  assign lines_5_ways_0_ready = (lines_5_ways_0_triggers[9 : 0] == 10'h000);
  assign io_contexts_10_staticWake = lines_5_ways_0_context_staticWake;
  assign io_contexts_10_physRd = lines_5_ways_0_context_physRd;
  assign io_contexts_10_robId = lines_5_ways_0_context_robId;
  assign io_contexts_10_euCtx_0 = lines_5_ways_0_context_euCtx_0;
  assign io_contexts_10_euCtx_1 = lines_5_ways_0_context_euCtx_1;
  always @(*) begin
    lines_5_ways_1_selComb = lines_5_ways_1_sel;
    if(lines_5_ways_1_fire) begin
      lines_5_ways_1_selComb = 2'b00;
    end
  end

  assign lines_5_ways_1_ready = (lines_5_ways_1_triggers[10 : 0] == 11'h000);
  assign io_contexts_11_staticWake = lines_5_ways_1_context_staticWake;
  assign io_contexts_11_physRd = lines_5_ways_1_context_physRd;
  assign io_contexts_11_robId = lines_5_ways_1_context_robId;
  assign io_contexts_11_euCtx_0 = lines_5_ways_1_context_euCtx_0;
  assign io_contexts_11_euCtx_1 = lines_5_ways_1_context_euCtx_1;
  always @(*) begin
    lines_6_ways_0_selComb = lines_6_ways_0_sel;
    if(lines_6_ways_0_fire) begin
      lines_6_ways_0_selComb = 2'b00;
    end
  end

  assign lines_6_ways_0_ready = (lines_6_ways_0_triggers[11 : 0] == 12'h000);
  assign io_contexts_12_staticWake = lines_6_ways_0_context_staticWake;
  assign io_contexts_12_physRd = lines_6_ways_0_context_physRd;
  assign io_contexts_12_robId = lines_6_ways_0_context_robId;
  assign io_contexts_12_euCtx_0 = lines_6_ways_0_context_euCtx_0;
  assign io_contexts_12_euCtx_1 = lines_6_ways_0_context_euCtx_1;
  always @(*) begin
    lines_6_ways_1_selComb = lines_6_ways_1_sel;
    if(lines_6_ways_1_fire) begin
      lines_6_ways_1_selComb = 2'b00;
    end
  end

  assign lines_6_ways_1_ready = (lines_6_ways_1_triggers[12 : 0] == 13'h0000);
  assign io_contexts_13_staticWake = lines_6_ways_1_context_staticWake;
  assign io_contexts_13_physRd = lines_6_ways_1_context_physRd;
  assign io_contexts_13_robId = lines_6_ways_1_context_robId;
  assign io_contexts_13_euCtx_0 = lines_6_ways_1_context_euCtx_0;
  assign io_contexts_13_euCtx_1 = lines_6_ways_1_context_euCtx_1;
  always @(*) begin
    lines_7_ways_0_selComb = lines_7_ways_0_sel;
    if(lines_7_ways_0_fire) begin
      lines_7_ways_0_selComb = 2'b00;
    end
  end

  assign lines_7_ways_0_ready = (lines_7_ways_0_triggers[13 : 0] == 14'h0000);
  assign io_contexts_14_staticWake = lines_7_ways_0_context_staticWake;
  assign io_contexts_14_physRd = lines_7_ways_0_context_physRd;
  assign io_contexts_14_robId = lines_7_ways_0_context_robId;
  assign io_contexts_14_euCtx_0 = lines_7_ways_0_context_euCtx_0;
  assign io_contexts_14_euCtx_1 = lines_7_ways_0_context_euCtx_1;
  always @(*) begin
    lines_7_ways_1_selComb = lines_7_ways_1_sel;
    if(lines_7_ways_1_fire) begin
      lines_7_ways_1_selComb = 2'b00;
    end
  end

  assign lines_7_ways_1_ready = (lines_7_ways_1_triggers[14 : 0] == 15'h0000);
  assign io_contexts_15_staticWake = lines_7_ways_1_context_staticWake;
  assign io_contexts_15_physRd = lines_7_ways_1_context_physRd;
  assign io_contexts_15_robId = lines_7_ways_1_context_robId;
  assign io_contexts_15_euCtx_0 = lines_7_ways_1_context_euCtx_0;
  assign io_contexts_15_euCtx_1 = lines_7_ways_1_context_euCtx_1;
  always @(*) begin
    lines_8_ways_0_selComb = lines_8_ways_0_sel;
    if(lines_8_ways_0_fire) begin
      lines_8_ways_0_selComb = 2'b00;
    end
  end

  assign lines_8_ways_0_ready = (lines_8_ways_0_triggers[15 : 0] == 16'h0000);
  assign io_contexts_16_staticWake = lines_8_ways_0_context_staticWake;
  assign io_contexts_16_physRd = lines_8_ways_0_context_physRd;
  assign io_contexts_16_robId = lines_8_ways_0_context_robId;
  assign io_contexts_16_euCtx_0 = lines_8_ways_0_context_euCtx_0;
  assign io_contexts_16_euCtx_1 = lines_8_ways_0_context_euCtx_1;
  always @(*) begin
    lines_8_ways_1_selComb = lines_8_ways_1_sel;
    if(lines_8_ways_1_fire) begin
      lines_8_ways_1_selComb = 2'b00;
    end
  end

  assign lines_8_ways_1_ready = (lines_8_ways_1_triggers[16 : 0] == 17'h00000);
  assign io_contexts_17_staticWake = lines_8_ways_1_context_staticWake;
  assign io_contexts_17_physRd = lines_8_ways_1_context_physRd;
  assign io_contexts_17_robId = lines_8_ways_1_context_robId;
  assign io_contexts_17_euCtx_0 = lines_8_ways_1_context_euCtx_0;
  assign io_contexts_17_euCtx_1 = lines_8_ways_1_context_euCtx_1;
  always @(*) begin
    lines_9_ways_0_selComb = lines_9_ways_0_sel;
    if(lines_9_ways_0_fire) begin
      lines_9_ways_0_selComb = 2'b00;
    end
  end

  assign lines_9_ways_0_ready = (lines_9_ways_0_triggers[17 : 0] == 18'h00000);
  assign io_contexts_18_staticWake = lines_9_ways_0_context_staticWake;
  assign io_contexts_18_physRd = lines_9_ways_0_context_physRd;
  assign io_contexts_18_robId = lines_9_ways_0_context_robId;
  assign io_contexts_18_euCtx_0 = lines_9_ways_0_context_euCtx_0;
  assign io_contexts_18_euCtx_1 = lines_9_ways_0_context_euCtx_1;
  always @(*) begin
    lines_9_ways_1_selComb = lines_9_ways_1_sel;
    if(lines_9_ways_1_fire) begin
      lines_9_ways_1_selComb = 2'b00;
    end
  end

  assign lines_9_ways_1_ready = (lines_9_ways_1_triggers[18 : 0] == 19'h00000);
  assign io_contexts_19_staticWake = lines_9_ways_1_context_staticWake;
  assign io_contexts_19_physRd = lines_9_ways_1_context_physRd;
  assign io_contexts_19_robId = lines_9_ways_1_context_robId;
  assign io_contexts_19_euCtx_0 = lines_9_ways_1_context_euCtx_0;
  assign io_contexts_19_euCtx_1 = lines_9_ways_1_context_euCtx_1;
  always @(*) begin
    lines_10_ways_0_selComb = lines_10_ways_0_sel;
    if(lines_10_ways_0_fire) begin
      lines_10_ways_0_selComb = 2'b00;
    end
  end

  assign lines_10_ways_0_ready = (lines_10_ways_0_triggers[19 : 0] == 20'h00000);
  assign io_contexts_20_staticWake = lines_10_ways_0_context_staticWake;
  assign io_contexts_20_physRd = lines_10_ways_0_context_physRd;
  assign io_contexts_20_robId = lines_10_ways_0_context_robId;
  assign io_contexts_20_euCtx_0 = lines_10_ways_0_context_euCtx_0;
  assign io_contexts_20_euCtx_1 = lines_10_ways_0_context_euCtx_1;
  always @(*) begin
    lines_10_ways_1_selComb = lines_10_ways_1_sel;
    if(lines_10_ways_1_fire) begin
      lines_10_ways_1_selComb = 2'b00;
    end
  end

  assign lines_10_ways_1_ready = (lines_10_ways_1_triggers[20 : 0] == 21'h000000);
  assign io_contexts_21_staticWake = lines_10_ways_1_context_staticWake;
  assign io_contexts_21_physRd = lines_10_ways_1_context_physRd;
  assign io_contexts_21_robId = lines_10_ways_1_context_robId;
  assign io_contexts_21_euCtx_0 = lines_10_ways_1_context_euCtx_0;
  assign io_contexts_21_euCtx_1 = lines_10_ways_1_context_euCtx_1;
  always @(*) begin
    lines_11_ways_0_selComb = lines_11_ways_0_sel;
    if(lines_11_ways_0_fire) begin
      lines_11_ways_0_selComb = 2'b00;
    end
  end

  assign lines_11_ways_0_ready = (lines_11_ways_0_triggers[21 : 0] == 22'h000000);
  assign io_contexts_22_staticWake = lines_11_ways_0_context_staticWake;
  assign io_contexts_22_physRd = lines_11_ways_0_context_physRd;
  assign io_contexts_22_robId = lines_11_ways_0_context_robId;
  assign io_contexts_22_euCtx_0 = lines_11_ways_0_context_euCtx_0;
  assign io_contexts_22_euCtx_1 = lines_11_ways_0_context_euCtx_1;
  always @(*) begin
    lines_11_ways_1_selComb = lines_11_ways_1_sel;
    if(lines_11_ways_1_fire) begin
      lines_11_ways_1_selComb = 2'b00;
    end
  end

  assign lines_11_ways_1_ready = (lines_11_ways_1_triggers[22 : 0] == 23'h000000);
  assign io_contexts_23_staticWake = lines_11_ways_1_context_staticWake;
  assign io_contexts_23_physRd = lines_11_ways_1_context_physRd;
  assign io_contexts_23_robId = lines_11_ways_1_context_robId;
  assign io_contexts_23_euCtx_0 = lines_11_ways_1_context_euCtx_0;
  assign io_contexts_23_euCtx_1 = lines_11_ways_1_context_euCtx_1;
  always @(*) begin
    lines_12_ways_0_selComb = lines_12_ways_0_sel;
    if(lines_12_ways_0_fire) begin
      lines_12_ways_0_selComb = 2'b00;
    end
  end

  assign lines_12_ways_0_ready = (lines_12_ways_0_triggers[23 : 0] == 24'h000000);
  assign io_contexts_24_staticWake = lines_12_ways_0_context_staticWake;
  assign io_contexts_24_physRd = lines_12_ways_0_context_physRd;
  assign io_contexts_24_robId = lines_12_ways_0_context_robId;
  assign io_contexts_24_euCtx_0 = lines_12_ways_0_context_euCtx_0;
  assign io_contexts_24_euCtx_1 = lines_12_ways_0_context_euCtx_1;
  always @(*) begin
    lines_12_ways_1_selComb = lines_12_ways_1_sel;
    if(lines_12_ways_1_fire) begin
      lines_12_ways_1_selComb = 2'b00;
    end
  end

  assign lines_12_ways_1_ready = (lines_12_ways_1_triggers[24 : 0] == 25'h0000000);
  assign io_contexts_25_staticWake = lines_12_ways_1_context_staticWake;
  assign io_contexts_25_physRd = lines_12_ways_1_context_physRd;
  assign io_contexts_25_robId = lines_12_ways_1_context_robId;
  assign io_contexts_25_euCtx_0 = lines_12_ways_1_context_euCtx_0;
  assign io_contexts_25_euCtx_1 = lines_12_ways_1_context_euCtx_1;
  always @(*) begin
    lines_13_ways_0_selComb = lines_13_ways_0_sel;
    if(lines_13_ways_0_fire) begin
      lines_13_ways_0_selComb = 2'b00;
    end
  end

  assign lines_13_ways_0_ready = (lines_13_ways_0_triggers[25 : 0] == 26'h0000000);
  assign io_contexts_26_staticWake = lines_13_ways_0_context_staticWake;
  assign io_contexts_26_physRd = lines_13_ways_0_context_physRd;
  assign io_contexts_26_robId = lines_13_ways_0_context_robId;
  assign io_contexts_26_euCtx_0 = lines_13_ways_0_context_euCtx_0;
  assign io_contexts_26_euCtx_1 = lines_13_ways_0_context_euCtx_1;
  always @(*) begin
    lines_13_ways_1_selComb = lines_13_ways_1_sel;
    if(lines_13_ways_1_fire) begin
      lines_13_ways_1_selComb = 2'b00;
    end
  end

  assign lines_13_ways_1_ready = (lines_13_ways_1_triggers[26 : 0] == 27'h0000000);
  assign io_contexts_27_staticWake = lines_13_ways_1_context_staticWake;
  assign io_contexts_27_physRd = lines_13_ways_1_context_physRd;
  assign io_contexts_27_robId = lines_13_ways_1_context_robId;
  assign io_contexts_27_euCtx_0 = lines_13_ways_1_context_euCtx_0;
  assign io_contexts_27_euCtx_1 = lines_13_ways_1_context_euCtx_1;
  always @(*) begin
    lines_14_ways_0_selComb = lines_14_ways_0_sel;
    if(lines_14_ways_0_fire) begin
      lines_14_ways_0_selComb = 2'b00;
    end
  end

  assign lines_14_ways_0_ready = (lines_14_ways_0_triggers[27 : 0] == 28'h0000000);
  assign io_contexts_28_staticWake = lines_14_ways_0_context_staticWake;
  assign io_contexts_28_physRd = lines_14_ways_0_context_physRd;
  assign io_contexts_28_robId = lines_14_ways_0_context_robId;
  assign io_contexts_28_euCtx_0 = lines_14_ways_0_context_euCtx_0;
  assign io_contexts_28_euCtx_1 = lines_14_ways_0_context_euCtx_1;
  always @(*) begin
    lines_14_ways_1_selComb = lines_14_ways_1_sel;
    if(lines_14_ways_1_fire) begin
      lines_14_ways_1_selComb = 2'b00;
    end
  end

  assign lines_14_ways_1_ready = (lines_14_ways_1_triggers[28 : 0] == 29'h00000000);
  assign io_contexts_29_staticWake = lines_14_ways_1_context_staticWake;
  assign io_contexts_29_physRd = lines_14_ways_1_context_physRd;
  assign io_contexts_29_robId = lines_14_ways_1_context_robId;
  assign io_contexts_29_euCtx_0 = lines_14_ways_1_context_euCtx_0;
  assign io_contexts_29_euCtx_1 = lines_14_ways_1_context_euCtx_1;
  always @(*) begin
    lines_15_ways_0_selComb = lines_15_ways_0_sel;
    if(lines_15_ways_0_fire) begin
      lines_15_ways_0_selComb = 2'b00;
    end
  end

  assign lines_15_ways_0_ready = (lines_15_ways_0_triggers[29 : 0] == 30'h00000000);
  assign io_contexts_30_staticWake = lines_15_ways_0_context_staticWake;
  assign io_contexts_30_physRd = lines_15_ways_0_context_physRd;
  assign io_contexts_30_robId = lines_15_ways_0_context_robId;
  assign io_contexts_30_euCtx_0 = lines_15_ways_0_context_euCtx_0;
  assign io_contexts_30_euCtx_1 = lines_15_ways_0_context_euCtx_1;
  always @(*) begin
    lines_15_ways_1_selComb = lines_15_ways_1_sel;
    if(lines_15_ways_1_fire) begin
      lines_15_ways_1_selComb = 2'b00;
    end
  end

  assign lines_15_ways_1_ready = (lines_15_ways_1_triggers[30 : 0] == 31'h00000000);
  assign io_contexts_31_staticWake = lines_15_ways_1_context_staticWake;
  assign io_contexts_31_physRd = lines_15_ways_1_context_physRd;
  assign io_contexts_31_robId = lines_15_ways_1_context_robId;
  assign io_contexts_31_euCtx_0 = lines_15_ways_1_context_euCtx_0;
  assign io_contexts_31_euCtx_1 = lines_15_ways_1_context_euCtx_1;
  assign compaction_moveIt = (io_push_valid && io_push_ready);
  assign event_moved = ((! compaction_moveIt) ? io_events : _zz_event_moved);
  assign event_value = (clear ? 32'hffffffff : event_moved);
  assign when_IssueQueue_l109 = event_value[0];
  assign when_IssueQueue_l109_1 = event_value[1];
  assign when_IssueQueue_l109_2 = event_value[2];
  assign when_IssueQueue_l109_3 = event_value[3];
  assign when_IssueQueue_l109_4 = event_value[4];
  assign when_IssueQueue_l109_5 = event_value[5];
  assign when_IssueQueue_l109_6 = event_value[6];
  assign when_IssueQueue_l109_7 = event_value[7];
  assign when_IssueQueue_l109_8 = event_value[8];
  assign when_IssueQueue_l109_9 = event_value[9];
  assign when_IssueQueue_l109_10 = event_value[10];
  assign when_IssueQueue_l109_11 = event_value[11];
  assign when_IssueQueue_l109_12 = event_value[12];
  assign when_IssueQueue_l109_13 = event_value[13];
  assign when_IssueQueue_l109_14 = event_value[14];
  assign when_IssueQueue_l109_15 = event_value[15];
  assign when_IssueQueue_l109_16 = event_value[16];
  assign when_IssueQueue_l109_17 = event_value[17];
  assign when_IssueQueue_l109_18 = event_value[18];
  assign when_IssueQueue_l109_19 = event_value[19];
  assign when_IssueQueue_l109_20 = event_value[20];
  assign when_IssueQueue_l109_21 = event_value[21];
  assign when_IssueQueue_l109_22 = event_value[22];
  assign when_IssueQueue_l109_23 = event_value[23];
  assign when_IssueQueue_l109_24 = event_value[24];
  assign when_IssueQueue_l109_25 = event_value[25];
  assign when_IssueQueue_l109_26 = event_value[26];
  assign when_IssueQueue_l109_27 = event_value[27];
  assign when_IssueQueue_l109_28 = event_value[28];
  assign when_IssueQueue_l109_29 = event_value[29];
  assign when_IssueQueue_l109_30 = event_value[30];
  assign when_IssueQueue_l109_31 = event_value[31];
  assign selector_0_slotsValid = {(lines_15_ways_0_ready && lines_15_ways_0_sel[0]),{(lines_14_ways_0_ready && lines_14_ways_0_sel[0]),{(lines_13_ways_0_ready && lines_13_ways_0_sel[0]),{(lines_12_ways_0_ready && lines_12_ways_0_sel[0]),{(lines_11_ways_0_ready && _zz_selector_0_slotsValid),{_zz_selector_0_slotsValid_1,{_zz_selector_0_slotsValid_2,_zz_selector_0_slotsValid_3}}}}}}};
  assign _zz_selector_0_slotsValid_bools_0 = selector_0_slotsValid;
  assign selector_0_slotsValid_bools_0 = _zz_selector_0_slotsValid_bools_0[0];
  assign selector_0_slotsValid_bools_1 = _zz_selector_0_slotsValid_bools_0[1];
  assign selector_0_slotsValid_bools_2 = _zz_selector_0_slotsValid_bools_0[2];
  assign selector_0_slotsValid_bools_3 = _zz_selector_0_slotsValid_bools_0[3];
  assign selector_0_slotsValid_bools_4 = _zz_selector_0_slotsValid_bools_0[4];
  assign selector_0_slotsValid_bools_5 = _zz_selector_0_slotsValid_bools_0[5];
  assign selector_0_slotsValid_bools_6 = _zz_selector_0_slotsValid_bools_0[6];
  assign selector_0_slotsValid_bools_7 = _zz_selector_0_slotsValid_bools_0[7];
  assign selector_0_slotsValid_bools_8 = _zz_selector_0_slotsValid_bools_0[8];
  assign selector_0_slotsValid_bools_9 = _zz_selector_0_slotsValid_bools_0[9];
  assign selector_0_slotsValid_bools_10 = _zz_selector_0_slotsValid_bools_0[10];
  assign selector_0_slotsValid_bools_11 = _zz_selector_0_slotsValid_bools_0[11];
  assign selector_0_slotsValid_bools_12 = _zz_selector_0_slotsValid_bools_0[12];
  assign selector_0_slotsValid_bools_13 = _zz_selector_0_slotsValid_bools_0[13];
  assign selector_0_slotsValid_bools_14 = _zz_selector_0_slotsValid_bools_0[14];
  assign selector_0_slotsValid_bools_15 = _zz_selector_0_slotsValid_bools_0[15];
  always @(*) begin
    _zz_selector_0_selOh[0] = (selector_0_slotsValid_bools_0 && (! 1'b0));
    _zz_selector_0_selOh[1] = (selector_0_slotsValid_bools_1 && (! selector_0_slotsValid_bools_0));
    _zz_selector_0_selOh[2] = (selector_0_slotsValid_bools_2 && (! selector_0_slotsValid_range_0_to_1));
    _zz_selector_0_selOh[3] = (selector_0_slotsValid_bools_3 && (! selector_0_slotsValid_range_0_to_2));
    _zz_selector_0_selOh[4] = (selector_0_slotsValid_bools_4 && (! selector_0_slotsValid_range_0_to_3));
    _zz_selector_0_selOh[5] = (selector_0_slotsValid_bools_5 && (! selector_0_slotsValid_range_0_to_4));
    _zz_selector_0_selOh[6] = (selector_0_slotsValid_bools_6 && (! selector_0_slotsValid_range_0_to_5));
    _zz_selector_0_selOh[7] = (selector_0_slotsValid_bools_7 && (! (selector_0_slotsValid_bools_6 || selector_0_slotsValid_range_0_to_5)));
    _zz_selector_0_selOh[8] = (selector_0_slotsValid_bools_8 && (! (selector_0_slotsValid_range_6_to_7 || selector_0_slotsValid_range_0_to_5)));
    _zz_selector_0_selOh[9] = (selector_0_slotsValid_bools_9 && (! (selector_0_slotsValid_range_6_to_8 || selector_0_slotsValid_range_0_to_5)));
    _zz_selector_0_selOh[10] = (selector_0_slotsValid_bools_10 && (! (selector_0_slotsValid_range_6_to_9 || selector_0_slotsValid_range_0_to_5)));
    _zz_selector_0_selOh[11] = (selector_0_slotsValid_bools_11 && (! (selector_0_slotsValid_range_6_to_10 || selector_0_slotsValid_range_0_to_5)));
    _zz_selector_0_selOh[12] = (selector_0_slotsValid_bools_12 && (! (selector_0_slotsValid_range_6_to_11 || selector_0_slotsValid_range_0_to_5)));
    _zz_selector_0_selOh[13] = (selector_0_slotsValid_bools_13 && (! (selector_0_slotsValid_bools_12 || selector_0_slotsValid_range_0_to_11)));
    _zz_selector_0_selOh[14] = (selector_0_slotsValid_bools_14 && (! (selector_0_slotsValid_range_12_to_13 || selector_0_slotsValid_range_0_to_11)));
    _zz_selector_0_selOh[15] = (selector_0_slotsValid_bools_15 && (! (selector_0_slotsValid_range_12_to_14 || selector_0_slotsValid_range_0_to_11)));
  end

  assign selector_0_slotsValid_range_0_to_1 = ({selector_0_slotsValid_bools_1,selector_0_slotsValid_bools_0} != 2'b00);
  assign selector_0_slotsValid_range_0_to_2 = ({selector_0_slotsValid_bools_2,{selector_0_slotsValid_bools_1,selector_0_slotsValid_bools_0}} != 3'b000);
  assign selector_0_slotsValid_range_0_to_3 = ({selector_0_slotsValid_bools_3,{selector_0_slotsValid_bools_2,{selector_0_slotsValid_bools_1,selector_0_slotsValid_bools_0}}} != 4'b0000);
  assign selector_0_slotsValid_range_0_to_4 = ({selector_0_slotsValid_bools_4,{selector_0_slotsValid_bools_3,{selector_0_slotsValid_bools_2,{selector_0_slotsValid_bools_1,selector_0_slotsValid_bools_0}}}} != 5'h00);
  assign selector_0_slotsValid_range_0_to_5 = ({selector_0_slotsValid_bools_5,{selector_0_slotsValid_bools_4,{selector_0_slotsValid_bools_3,{selector_0_slotsValid_bools_2,{selector_0_slotsValid_bools_1,selector_0_slotsValid_bools_0}}}}} != 6'h00);
  assign selector_0_slotsValid_range_6_to_7 = ({selector_0_slotsValid_bools_7,selector_0_slotsValid_bools_6} != 2'b00);
  assign selector_0_slotsValid_range_6_to_8 = ({selector_0_slotsValid_bools_8,{selector_0_slotsValid_bools_7,selector_0_slotsValid_bools_6}} != 3'b000);
  assign selector_0_slotsValid_range_6_to_9 = ({selector_0_slotsValid_bools_9,{selector_0_slotsValid_bools_8,{selector_0_slotsValid_bools_7,selector_0_slotsValid_bools_6}}} != 4'b0000);
  assign selector_0_slotsValid_range_6_to_10 = ({selector_0_slotsValid_bools_10,{selector_0_slotsValid_bools_9,{selector_0_slotsValid_bools_8,{selector_0_slotsValid_bools_7,selector_0_slotsValid_bools_6}}}} != 5'h00);
  assign selector_0_slotsValid_range_6_to_11 = ({selector_0_slotsValid_bools_11,{selector_0_slotsValid_bools_10,{selector_0_slotsValid_bools_9,{selector_0_slotsValid_bools_8,{selector_0_slotsValid_bools_7,selector_0_slotsValid_bools_6}}}}} != 6'h00);
  assign selector_0_slotsValid_range_0_to_11 = ({selector_0_slotsValid_range_6_to_11,selector_0_slotsValid_range_0_to_5} != 2'b00);
  assign selector_0_slotsValid_range_12_to_13 = ({selector_0_slotsValid_bools_13,selector_0_slotsValid_bools_12} != 2'b00);
  assign selector_0_slotsValid_range_12_to_14 = ({selector_0_slotsValid_bools_14,{selector_0_slotsValid_bools_13,selector_0_slotsValid_bools_12}} != 3'b000);
  assign selector_0_selOh = _zz_selector_0_selOh;
  assign io_schedules_0_valid = ((|selector_0_slotsValid) && running);
  assign io_schedules_0_payload_event = selector_0_selOh;
  assign selector_1_slotsValid = {(lines_15_ways_1_ready && lines_15_ways_1_sel[0]),{(lines_14_ways_1_ready && lines_14_ways_1_sel[0]),{(lines_13_ways_1_ready && lines_13_ways_1_sel[0]),{(lines_12_ways_1_ready && lines_12_ways_1_sel[0]),{(lines_11_ways_1_ready && _zz_selector_1_slotsValid),{_zz_selector_1_slotsValid_1,{_zz_selector_1_slotsValid_2,_zz_selector_1_slotsValid_3}}}}}}};
  assign _zz_selector_1_slotsValid_bools_0 = selector_1_slotsValid;
  assign selector_1_slotsValid_bools_0 = _zz_selector_1_slotsValid_bools_0[0];
  assign selector_1_slotsValid_bools_1 = _zz_selector_1_slotsValid_bools_0[1];
  assign selector_1_slotsValid_bools_2 = _zz_selector_1_slotsValid_bools_0[2];
  assign selector_1_slotsValid_bools_3 = _zz_selector_1_slotsValid_bools_0[3];
  assign selector_1_slotsValid_bools_4 = _zz_selector_1_slotsValid_bools_0[4];
  assign selector_1_slotsValid_bools_5 = _zz_selector_1_slotsValid_bools_0[5];
  assign selector_1_slotsValid_bools_6 = _zz_selector_1_slotsValid_bools_0[6];
  assign selector_1_slotsValid_bools_7 = _zz_selector_1_slotsValid_bools_0[7];
  assign selector_1_slotsValid_bools_8 = _zz_selector_1_slotsValid_bools_0[8];
  assign selector_1_slotsValid_bools_9 = _zz_selector_1_slotsValid_bools_0[9];
  assign selector_1_slotsValid_bools_10 = _zz_selector_1_slotsValid_bools_0[10];
  assign selector_1_slotsValid_bools_11 = _zz_selector_1_slotsValid_bools_0[11];
  assign selector_1_slotsValid_bools_12 = _zz_selector_1_slotsValid_bools_0[12];
  assign selector_1_slotsValid_bools_13 = _zz_selector_1_slotsValid_bools_0[13];
  assign selector_1_slotsValid_bools_14 = _zz_selector_1_slotsValid_bools_0[14];
  assign selector_1_slotsValid_bools_15 = _zz_selector_1_slotsValid_bools_0[15];
  always @(*) begin
    _zz_selector_1_selOh[0] = (selector_1_slotsValid_bools_0 && (! 1'b0));
    _zz_selector_1_selOh[1] = (selector_1_slotsValid_bools_1 && (! selector_1_slotsValid_bools_0));
    _zz_selector_1_selOh[2] = (selector_1_slotsValid_bools_2 && (! selector_1_slotsValid_range_0_to_1));
    _zz_selector_1_selOh[3] = (selector_1_slotsValid_bools_3 && (! selector_1_slotsValid_range_0_to_2));
    _zz_selector_1_selOh[4] = (selector_1_slotsValid_bools_4 && (! selector_1_slotsValid_range_0_to_3));
    _zz_selector_1_selOh[5] = (selector_1_slotsValid_bools_5 && (! selector_1_slotsValid_range_0_to_4));
    _zz_selector_1_selOh[6] = (selector_1_slotsValid_bools_6 && (! selector_1_slotsValid_range_0_to_5));
    _zz_selector_1_selOh[7] = (selector_1_slotsValid_bools_7 && (! (selector_1_slotsValid_bools_6 || selector_1_slotsValid_range_0_to_5)));
    _zz_selector_1_selOh[8] = (selector_1_slotsValid_bools_8 && (! (selector_1_slotsValid_range_6_to_7 || selector_1_slotsValid_range_0_to_5)));
    _zz_selector_1_selOh[9] = (selector_1_slotsValid_bools_9 && (! (selector_1_slotsValid_range_6_to_8 || selector_1_slotsValid_range_0_to_5)));
    _zz_selector_1_selOh[10] = (selector_1_slotsValid_bools_10 && (! (selector_1_slotsValid_range_6_to_9 || selector_1_slotsValid_range_0_to_5)));
    _zz_selector_1_selOh[11] = (selector_1_slotsValid_bools_11 && (! (selector_1_slotsValid_range_6_to_10 || selector_1_slotsValid_range_0_to_5)));
    _zz_selector_1_selOh[12] = (selector_1_slotsValid_bools_12 && (! (selector_1_slotsValid_range_6_to_11 || selector_1_slotsValid_range_0_to_5)));
    _zz_selector_1_selOh[13] = (selector_1_slotsValid_bools_13 && (! (selector_1_slotsValid_bools_12 || selector_1_slotsValid_range_0_to_11)));
    _zz_selector_1_selOh[14] = (selector_1_slotsValid_bools_14 && (! (selector_1_slotsValid_range_12_to_13 || selector_1_slotsValid_range_0_to_11)));
    _zz_selector_1_selOh[15] = (selector_1_slotsValid_bools_15 && (! (selector_1_slotsValid_range_12_to_14 || selector_1_slotsValid_range_0_to_11)));
  end

  assign selector_1_slotsValid_range_0_to_1 = ({selector_1_slotsValid_bools_1,selector_1_slotsValid_bools_0} != 2'b00);
  assign selector_1_slotsValid_range_0_to_2 = ({selector_1_slotsValid_bools_2,{selector_1_slotsValid_bools_1,selector_1_slotsValid_bools_0}} != 3'b000);
  assign selector_1_slotsValid_range_0_to_3 = ({selector_1_slotsValid_bools_3,{selector_1_slotsValid_bools_2,{selector_1_slotsValid_bools_1,selector_1_slotsValid_bools_0}}} != 4'b0000);
  assign selector_1_slotsValid_range_0_to_4 = ({selector_1_slotsValid_bools_4,{selector_1_slotsValid_bools_3,{selector_1_slotsValid_bools_2,{selector_1_slotsValid_bools_1,selector_1_slotsValid_bools_0}}}} != 5'h00);
  assign selector_1_slotsValid_range_0_to_5 = ({selector_1_slotsValid_bools_5,{selector_1_slotsValid_bools_4,{selector_1_slotsValid_bools_3,{selector_1_slotsValid_bools_2,{selector_1_slotsValid_bools_1,selector_1_slotsValid_bools_0}}}}} != 6'h00);
  assign selector_1_slotsValid_range_6_to_7 = ({selector_1_slotsValid_bools_7,selector_1_slotsValid_bools_6} != 2'b00);
  assign selector_1_slotsValid_range_6_to_8 = ({selector_1_slotsValid_bools_8,{selector_1_slotsValid_bools_7,selector_1_slotsValid_bools_6}} != 3'b000);
  assign selector_1_slotsValid_range_6_to_9 = ({selector_1_slotsValid_bools_9,{selector_1_slotsValid_bools_8,{selector_1_slotsValid_bools_7,selector_1_slotsValid_bools_6}}} != 4'b0000);
  assign selector_1_slotsValid_range_6_to_10 = ({selector_1_slotsValid_bools_10,{selector_1_slotsValid_bools_9,{selector_1_slotsValid_bools_8,{selector_1_slotsValid_bools_7,selector_1_slotsValid_bools_6}}}} != 5'h00);
  assign selector_1_slotsValid_range_6_to_11 = ({selector_1_slotsValid_bools_11,{selector_1_slotsValid_bools_10,{selector_1_slotsValid_bools_9,{selector_1_slotsValid_bools_8,{selector_1_slotsValid_bools_7,selector_1_slotsValid_bools_6}}}}} != 6'h00);
  assign selector_1_slotsValid_range_0_to_11 = ({selector_1_slotsValid_range_6_to_11,selector_1_slotsValid_range_0_to_5} != 2'b00);
  assign selector_1_slotsValid_range_12_to_13 = ({selector_1_slotsValid_bools_13,selector_1_slotsValid_bools_12} != 2'b00);
  assign selector_1_slotsValid_range_12_to_14 = ({selector_1_slotsValid_bools_14,{selector_1_slotsValid_bools_13,selector_1_slotsValid_bools_12}} != 3'b000);
  assign selector_1_selOh = _zz_selector_1_selOh;
  assign io_schedules_1_valid = ((|selector_1_slotsValid) && running);
  assign io_schedules_1_payload_event = selector_1_selOh;
  assign selector_2_slotsValid = {(lines_15_ways_1_ready && lines_15_ways_1_sel[1]),{(lines_15_ways_0_ready && lines_15_ways_0_sel[1]),{(lines_14_ways_1_ready && lines_14_ways_1_sel[1]),{(lines_14_ways_0_ready && lines_14_ways_0_sel[1]),{(lines_13_ways_1_ready && _zz_selector_2_slotsValid),{_zz_selector_2_slotsValid_1,{_zz_selector_2_slotsValid_2,_zz_selector_2_slotsValid_3}}}}}}};
  assign _zz_selector_2_slotsValid_bools_0 = selector_2_slotsValid;
  assign selector_2_slotsValid_bools_0 = _zz_selector_2_slotsValid_bools_0[0];
  assign selector_2_slotsValid_bools_1 = _zz_selector_2_slotsValid_bools_0[1];
  assign selector_2_slotsValid_bools_2 = _zz_selector_2_slotsValid_bools_0[2];
  assign selector_2_slotsValid_bools_3 = _zz_selector_2_slotsValid_bools_0[3];
  assign selector_2_slotsValid_bools_4 = _zz_selector_2_slotsValid_bools_0[4];
  assign selector_2_slotsValid_bools_5 = _zz_selector_2_slotsValid_bools_0[5];
  assign selector_2_slotsValid_bools_6 = _zz_selector_2_slotsValid_bools_0[6];
  assign selector_2_slotsValid_bools_7 = _zz_selector_2_slotsValid_bools_0[7];
  assign selector_2_slotsValid_bools_8 = _zz_selector_2_slotsValid_bools_0[8];
  assign selector_2_slotsValid_bools_9 = _zz_selector_2_slotsValid_bools_0[9];
  assign selector_2_slotsValid_bools_10 = _zz_selector_2_slotsValid_bools_0[10];
  assign selector_2_slotsValid_bools_11 = _zz_selector_2_slotsValid_bools_0[11];
  assign selector_2_slotsValid_bools_12 = _zz_selector_2_slotsValid_bools_0[12];
  assign selector_2_slotsValid_bools_13 = _zz_selector_2_slotsValid_bools_0[13];
  assign selector_2_slotsValid_bools_14 = _zz_selector_2_slotsValid_bools_0[14];
  assign selector_2_slotsValid_bools_15 = _zz_selector_2_slotsValid_bools_0[15];
  assign selector_2_slotsValid_bools_16 = _zz_selector_2_slotsValid_bools_0[16];
  assign selector_2_slotsValid_bools_17 = _zz_selector_2_slotsValid_bools_0[17];
  assign selector_2_slotsValid_bools_18 = _zz_selector_2_slotsValid_bools_0[18];
  assign selector_2_slotsValid_bools_19 = _zz_selector_2_slotsValid_bools_0[19];
  assign selector_2_slotsValid_bools_20 = _zz_selector_2_slotsValid_bools_0[20];
  assign selector_2_slotsValid_bools_21 = _zz_selector_2_slotsValid_bools_0[21];
  assign selector_2_slotsValid_bools_22 = _zz_selector_2_slotsValid_bools_0[22];
  assign selector_2_slotsValid_bools_23 = _zz_selector_2_slotsValid_bools_0[23];
  assign selector_2_slotsValid_bools_24 = _zz_selector_2_slotsValid_bools_0[24];
  assign selector_2_slotsValid_bools_25 = _zz_selector_2_slotsValid_bools_0[25];
  assign selector_2_slotsValid_bools_26 = _zz_selector_2_slotsValid_bools_0[26];
  assign selector_2_slotsValid_bools_27 = _zz_selector_2_slotsValid_bools_0[27];
  assign selector_2_slotsValid_bools_28 = _zz_selector_2_slotsValid_bools_0[28];
  assign selector_2_slotsValid_bools_29 = _zz_selector_2_slotsValid_bools_0[29];
  assign selector_2_slotsValid_bools_30 = _zz_selector_2_slotsValid_bools_0[30];
  assign selector_2_slotsValid_bools_31 = _zz_selector_2_slotsValid_bools_0[31];
  always @(*) begin
    _zz_selector_2_selOh[0] = (selector_2_slotsValid_bools_0 && (! 1'b0));
    _zz_selector_2_selOh[1] = (selector_2_slotsValid_bools_1 && (! selector_2_slotsValid_bools_0));
    _zz_selector_2_selOh[2] = (selector_2_slotsValid_bools_2 && (! selector_2_slotsValid_range_0_to_1));
    _zz_selector_2_selOh[3] = (selector_2_slotsValid_bools_3 && (! selector_2_slotsValid_range_0_to_2));
    _zz_selector_2_selOh[4] = (selector_2_slotsValid_bools_4 && (! selector_2_slotsValid_range_0_to_3));
    _zz_selector_2_selOh[5] = (selector_2_slotsValid_bools_5 && (! selector_2_slotsValid_range_0_to_4));
    _zz_selector_2_selOh[6] = (selector_2_slotsValid_bools_6 && (! selector_2_slotsValid_range_0_to_5));
    _zz_selector_2_selOh[7] = (selector_2_slotsValid_bools_7 && (! (selector_2_slotsValid_bools_6 || selector_2_slotsValid_range_0_to_5)));
    _zz_selector_2_selOh[8] = (selector_2_slotsValid_bools_8 && (! (selector_2_slotsValid_range_6_to_7 || selector_2_slotsValid_range_0_to_5)));
    _zz_selector_2_selOh[9] = (selector_2_slotsValid_bools_9 && (! (selector_2_slotsValid_range_6_to_8 || selector_2_slotsValid_range_0_to_5)));
    _zz_selector_2_selOh[10] = (selector_2_slotsValid_bools_10 && (! (selector_2_slotsValid_range_6_to_9 || selector_2_slotsValid_range_0_to_5)));
    _zz_selector_2_selOh[11] = (selector_2_slotsValid_bools_11 && (! (selector_2_slotsValid_range_6_to_10 || selector_2_slotsValid_range_0_to_5)));
    _zz_selector_2_selOh[12] = (selector_2_slotsValid_bools_12 && (! (selector_2_slotsValid_range_6_to_11 || selector_2_slotsValid_range_0_to_5)));
    _zz_selector_2_selOh[13] = (selector_2_slotsValid_bools_13 && (! (selector_2_slotsValid_bools_12 || selector_2_slotsValid_range_0_to_11)));
    _zz_selector_2_selOh[14] = (selector_2_slotsValid_bools_14 && (! (selector_2_slotsValid_range_12_to_13 || selector_2_slotsValid_range_0_to_11)));
    _zz_selector_2_selOh[15] = (selector_2_slotsValid_bools_15 && (! (selector_2_slotsValid_range_12_to_14 || selector_2_slotsValid_range_0_to_11)));
    _zz_selector_2_selOh[16] = (selector_2_slotsValid_bools_16 && (! (selector_2_slotsValid_range_12_to_15 || selector_2_slotsValid_range_0_to_11)));
    _zz_selector_2_selOh[17] = (selector_2_slotsValid_bools_17 && (! (selector_2_slotsValid_range_12_to_16 || selector_2_slotsValid_range_0_to_11)));
    _zz_selector_2_selOh[18] = (selector_2_slotsValid_bools_18 && (! (selector_2_slotsValid_range_12_to_17 || selector_2_slotsValid_range_0_to_11)));
    _zz_selector_2_selOh[19] = (selector_2_slotsValid_bools_19 && (! (selector_2_slotsValid_bools_18 || selector_2_slotsValid_range_0_to_17)));
    _zz_selector_2_selOh[20] = (selector_2_slotsValid_bools_20 && (! (selector_2_slotsValid_range_18_to_19 || selector_2_slotsValid_range_0_to_17)));
    _zz_selector_2_selOh[21] = (selector_2_slotsValid_bools_21 && (! (selector_2_slotsValid_range_18_to_20 || selector_2_slotsValid_range_0_to_17)));
    _zz_selector_2_selOh[22] = (selector_2_slotsValid_bools_22 && (! (selector_2_slotsValid_range_18_to_21 || selector_2_slotsValid_range_0_to_17)));
    _zz_selector_2_selOh[23] = (selector_2_slotsValid_bools_23 && (! (selector_2_slotsValid_range_18_to_22 || selector_2_slotsValid_range_0_to_17)));
    _zz_selector_2_selOh[24] = (selector_2_slotsValid_bools_24 && (! (selector_2_slotsValid_range_18_to_23 || selector_2_slotsValid_range_0_to_17)));
    _zz_selector_2_selOh[25] = (selector_2_slotsValid_bools_25 && (! (selector_2_slotsValid_bools_24 || selector_2_slotsValid_range_0_to_23)));
    _zz_selector_2_selOh[26] = (selector_2_slotsValid_bools_26 && (! (selector_2_slotsValid_range_24_to_25 || selector_2_slotsValid_range_0_to_23)));
    _zz_selector_2_selOh[27] = (selector_2_slotsValid_bools_27 && (! (selector_2_slotsValid_range_24_to_26 || selector_2_slotsValid_range_0_to_23)));
    _zz_selector_2_selOh[28] = (selector_2_slotsValid_bools_28 && (! (selector_2_slotsValid_range_24_to_27 || selector_2_slotsValid_range_0_to_23)));
    _zz_selector_2_selOh[29] = (selector_2_slotsValid_bools_29 && (! (selector_2_slotsValid_range_24_to_28 || selector_2_slotsValid_range_0_to_23)));
    _zz_selector_2_selOh[30] = (selector_2_slotsValid_bools_30 && (! (selector_2_slotsValid_range_24_to_29 || selector_2_slotsValid_range_0_to_23)));
    _zz_selector_2_selOh[31] = (selector_2_slotsValid_bools_31 && (! (selector_2_slotsValid_bools_30 || selector_2_slotsValid_range_0_to_29)));
  end

  assign selector_2_slotsValid_range_0_to_1 = ({selector_2_slotsValid_bools_1,selector_2_slotsValid_bools_0} != 2'b00);
  assign selector_2_slotsValid_range_0_to_2 = ({selector_2_slotsValid_bools_2,{selector_2_slotsValid_bools_1,selector_2_slotsValid_bools_0}} != 3'b000);
  assign selector_2_slotsValid_range_0_to_3 = ({selector_2_slotsValid_bools_3,{selector_2_slotsValid_bools_2,{selector_2_slotsValid_bools_1,selector_2_slotsValid_bools_0}}} != 4'b0000);
  assign selector_2_slotsValid_range_0_to_4 = ({selector_2_slotsValid_bools_4,{selector_2_slotsValid_bools_3,{selector_2_slotsValid_bools_2,{selector_2_slotsValid_bools_1,selector_2_slotsValid_bools_0}}}} != 5'h00);
  assign selector_2_slotsValid_range_0_to_5 = ({selector_2_slotsValid_bools_5,{selector_2_slotsValid_bools_4,{selector_2_slotsValid_bools_3,{selector_2_slotsValid_bools_2,{selector_2_slotsValid_bools_1,selector_2_slotsValid_bools_0}}}}} != 6'h00);
  assign selector_2_slotsValid_range_6_to_7 = ({selector_2_slotsValid_bools_7,selector_2_slotsValid_bools_6} != 2'b00);
  assign selector_2_slotsValid_range_6_to_8 = ({selector_2_slotsValid_bools_8,{selector_2_slotsValid_bools_7,selector_2_slotsValid_bools_6}} != 3'b000);
  assign selector_2_slotsValid_range_6_to_9 = ({selector_2_slotsValid_bools_9,{selector_2_slotsValid_bools_8,{selector_2_slotsValid_bools_7,selector_2_slotsValid_bools_6}}} != 4'b0000);
  assign selector_2_slotsValid_range_6_to_10 = ({selector_2_slotsValid_bools_10,{selector_2_slotsValid_bools_9,{selector_2_slotsValid_bools_8,{selector_2_slotsValid_bools_7,selector_2_slotsValid_bools_6}}}} != 5'h00);
  assign selector_2_slotsValid_range_6_to_11 = ({selector_2_slotsValid_bools_11,{selector_2_slotsValid_bools_10,{selector_2_slotsValid_bools_9,{selector_2_slotsValid_bools_8,{selector_2_slotsValid_bools_7,selector_2_slotsValid_bools_6}}}}} != 6'h00);
  assign selector_2_slotsValid_range_0_to_11 = ({selector_2_slotsValid_range_6_to_11,selector_2_slotsValid_range_0_to_5} != 2'b00);
  assign selector_2_slotsValid_range_12_to_13 = ({selector_2_slotsValid_bools_13,selector_2_slotsValid_bools_12} != 2'b00);
  assign selector_2_slotsValid_range_12_to_14 = ({selector_2_slotsValid_bools_14,{selector_2_slotsValid_bools_13,selector_2_slotsValid_bools_12}} != 3'b000);
  assign selector_2_slotsValid_range_12_to_15 = ({selector_2_slotsValid_bools_15,{selector_2_slotsValid_bools_14,{selector_2_slotsValid_bools_13,selector_2_slotsValid_bools_12}}} != 4'b0000);
  assign selector_2_slotsValid_range_12_to_16 = ({selector_2_slotsValid_bools_16,{selector_2_slotsValid_bools_15,{selector_2_slotsValid_bools_14,{selector_2_slotsValid_bools_13,selector_2_slotsValid_bools_12}}}} != 5'h00);
  assign selector_2_slotsValid_range_12_to_17 = ({selector_2_slotsValid_bools_17,{selector_2_slotsValid_bools_16,{selector_2_slotsValid_bools_15,{selector_2_slotsValid_bools_14,{selector_2_slotsValid_bools_13,selector_2_slotsValid_bools_12}}}}} != 6'h00);
  assign selector_2_slotsValid_range_0_to_17 = ({selector_2_slotsValid_range_12_to_17,{selector_2_slotsValid_range_6_to_11,selector_2_slotsValid_range_0_to_5}} != 3'b000);
  assign selector_2_slotsValid_range_18_to_19 = ({selector_2_slotsValid_bools_19,selector_2_slotsValid_bools_18} != 2'b00);
  assign selector_2_slotsValid_range_18_to_20 = ({selector_2_slotsValid_bools_20,{selector_2_slotsValid_bools_19,selector_2_slotsValid_bools_18}} != 3'b000);
  assign selector_2_slotsValid_range_18_to_21 = ({selector_2_slotsValid_bools_21,{selector_2_slotsValid_bools_20,{selector_2_slotsValid_bools_19,selector_2_slotsValid_bools_18}}} != 4'b0000);
  assign selector_2_slotsValid_range_18_to_22 = ({selector_2_slotsValid_bools_22,{selector_2_slotsValid_bools_21,{selector_2_slotsValid_bools_20,{selector_2_slotsValid_bools_19,selector_2_slotsValid_bools_18}}}} != 5'h00);
  assign selector_2_slotsValid_range_18_to_23 = ({selector_2_slotsValid_bools_23,{selector_2_slotsValid_bools_22,{selector_2_slotsValid_bools_21,{selector_2_slotsValid_bools_20,{selector_2_slotsValid_bools_19,selector_2_slotsValid_bools_18}}}}} != 6'h00);
  assign selector_2_slotsValid_range_0_to_23 = ({selector_2_slotsValid_range_18_to_23,{selector_2_slotsValid_range_12_to_17,{selector_2_slotsValid_range_6_to_11,selector_2_slotsValid_range_0_to_5}}} != 4'b0000);
  assign selector_2_slotsValid_range_24_to_25 = ({selector_2_slotsValid_bools_25,selector_2_slotsValid_bools_24} != 2'b00);
  assign selector_2_slotsValid_range_24_to_26 = ({selector_2_slotsValid_bools_26,{selector_2_slotsValid_bools_25,selector_2_slotsValid_bools_24}} != 3'b000);
  assign selector_2_slotsValid_range_24_to_27 = ({selector_2_slotsValid_bools_27,{selector_2_slotsValid_bools_26,{selector_2_slotsValid_bools_25,selector_2_slotsValid_bools_24}}} != 4'b0000);
  assign selector_2_slotsValid_range_24_to_28 = ({selector_2_slotsValid_bools_28,{selector_2_slotsValid_bools_27,{selector_2_slotsValid_bools_26,{selector_2_slotsValid_bools_25,selector_2_slotsValid_bools_24}}}} != 5'h00);
  assign selector_2_slotsValid_range_24_to_29 = ({selector_2_slotsValid_bools_29,{selector_2_slotsValid_bools_28,{selector_2_slotsValid_bools_27,{selector_2_slotsValid_bools_26,{selector_2_slotsValid_bools_25,selector_2_slotsValid_bools_24}}}}} != 6'h00);
  assign selector_2_slotsValid_range_0_to_29 = ({selector_2_slotsValid_range_24_to_29,{selector_2_slotsValid_range_18_to_23,{selector_2_slotsValid_range_12_to_17,{selector_2_slotsValid_range_6_to_11,selector_2_slotsValid_range_0_to_5}}}} != 5'h00);
  assign selector_2_selOh = _zz_selector_2_selOh;
  assign io_schedules_2_valid = ((|selector_2_slotsValid) && running);
  assign io_schedules_2_payload_event = selector_2_selOh;
  assign lines_0_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[0]),(io_schedules_0_ready && selector_0_selOh[0])} != 2'b00);
  assign lines_0_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[1]),(io_schedules_1_ready && selector_1_selOh[0])} != 2'b00);
  assign lines_1_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[2]),(io_schedules_0_ready && selector_0_selOh[1])} != 2'b00);
  assign lines_1_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[3]),(io_schedules_1_ready && selector_1_selOh[1])} != 2'b00);
  assign lines_2_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[4]),(io_schedules_0_ready && selector_0_selOh[2])} != 2'b00);
  assign lines_2_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[5]),(io_schedules_1_ready && selector_1_selOh[2])} != 2'b00);
  assign lines_3_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[6]),(io_schedules_0_ready && selector_0_selOh[3])} != 2'b00);
  assign lines_3_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[7]),(io_schedules_1_ready && selector_1_selOh[3])} != 2'b00);
  assign lines_4_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[8]),(io_schedules_0_ready && selector_0_selOh[4])} != 2'b00);
  assign lines_4_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[9]),(io_schedules_1_ready && selector_1_selOh[4])} != 2'b00);
  assign lines_5_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[10]),(io_schedules_0_ready && selector_0_selOh[5])} != 2'b00);
  assign lines_5_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[11]),(io_schedules_1_ready && selector_1_selOh[5])} != 2'b00);
  assign lines_6_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[12]),(io_schedules_0_ready && selector_0_selOh[6])} != 2'b00);
  assign lines_6_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[13]),(io_schedules_1_ready && selector_1_selOh[6])} != 2'b00);
  assign lines_7_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[14]),(io_schedules_0_ready && selector_0_selOh[7])} != 2'b00);
  assign lines_7_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[15]),(io_schedules_1_ready && selector_1_selOh[7])} != 2'b00);
  assign lines_8_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[16]),(io_schedules_0_ready && selector_0_selOh[8])} != 2'b00);
  assign lines_8_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[17]),(io_schedules_1_ready && selector_1_selOh[8])} != 2'b00);
  assign lines_9_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[18]),(io_schedules_0_ready && selector_0_selOh[9])} != 2'b00);
  assign lines_9_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[19]),(io_schedules_1_ready && selector_1_selOh[9])} != 2'b00);
  assign lines_10_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[20]),(io_schedules_0_ready && selector_0_selOh[10])} != 2'b00);
  assign lines_10_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[21]),(io_schedules_1_ready && selector_1_selOh[10])} != 2'b00);
  assign lines_11_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[22]),(io_schedules_0_ready && selector_0_selOh[11])} != 2'b00);
  assign lines_11_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[23]),(io_schedules_1_ready && selector_1_selOh[11])} != 2'b00);
  assign lines_12_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[24]),(io_schedules_0_ready && selector_0_selOh[12])} != 2'b00);
  assign lines_12_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[25]),(io_schedules_1_ready && selector_1_selOh[12])} != 2'b00);
  assign lines_13_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[26]),(io_schedules_0_ready && selector_0_selOh[13])} != 2'b00);
  assign lines_13_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[27]),(io_schedules_1_ready && selector_1_selOh[13])} != 2'b00);
  assign lines_14_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[28]),(io_schedules_0_ready && selector_0_selOh[14])} != 2'b00);
  assign lines_14_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[29]),(io_schedules_1_ready && selector_1_selOh[14])} != 2'b00);
  assign lines_15_ways_0_fire = ({(io_schedules_2_ready && selector_2_selOh[30]),(io_schedules_0_ready && selector_0_selOh[15])} != 2'b00);
  assign lines_15_ways_1_fire = ({(io_schedules_2_ready && selector_2_selOh[31]),(io_schedules_1_ready && selector_1_selOh[15])} != 2'b00);
  assign line0Ready = (((! lines_0_ways_0_triggers[0]) && (lines_0_ways_0_sel == 2'b00)) && ((! lines_0_ways_1_triggers[1]) && (lines_0_ways_1_sel == 2'b00)));
  assign line1Ready = (((! lines_1_ways_0_triggers[2]) && (lines_1_ways_0_sel == 2'b00)) && ((! lines_1_ways_1_triggers[3]) && (lines_1_ways_1_sel == 2'b00)));
  assign io_push_ready = readyReg;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      running <= 1'b0;
      readyReg <= 1'b0;
    end else begin
      running <= 1'b1;
      readyReg <= (compaction_moveIt ? line1Ready : line0Ready);
    end
  end

  always @(posedge clk) begin
    lines_0_ways_0_sel <= lines_0_ways_0_selComb;
    lines_0_ways_1_sel <= lines_0_ways_1_selComb;
    lines_1_ways_0_sel <= lines_1_ways_0_selComb;
    lines_1_ways_1_sel <= lines_1_ways_1_selComb;
    lines_2_ways_0_sel <= lines_2_ways_0_selComb;
    lines_2_ways_1_sel <= lines_2_ways_1_selComb;
    lines_3_ways_0_sel <= lines_3_ways_0_selComb;
    lines_3_ways_1_sel <= lines_3_ways_1_selComb;
    lines_4_ways_0_sel <= lines_4_ways_0_selComb;
    lines_4_ways_1_sel <= lines_4_ways_1_selComb;
    lines_5_ways_0_sel <= lines_5_ways_0_selComb;
    lines_5_ways_1_sel <= lines_5_ways_1_selComb;
    lines_6_ways_0_sel <= lines_6_ways_0_selComb;
    lines_6_ways_1_sel <= lines_6_ways_1_selComb;
    lines_7_ways_0_sel <= lines_7_ways_0_selComb;
    lines_7_ways_1_sel <= lines_7_ways_1_selComb;
    lines_8_ways_0_sel <= lines_8_ways_0_selComb;
    lines_8_ways_1_sel <= lines_8_ways_1_selComb;
    lines_9_ways_0_sel <= lines_9_ways_0_selComb;
    lines_9_ways_1_sel <= lines_9_ways_1_selComb;
    lines_10_ways_0_sel <= lines_10_ways_0_selComb;
    lines_10_ways_1_sel <= lines_10_ways_1_selComb;
    lines_11_ways_0_sel <= lines_11_ways_0_selComb;
    lines_11_ways_1_sel <= lines_11_ways_1_selComb;
    lines_12_ways_0_sel <= lines_12_ways_0_selComb;
    lines_12_ways_1_sel <= lines_12_ways_1_selComb;
    lines_13_ways_0_sel <= lines_13_ways_0_selComb;
    lines_13_ways_1_sel <= lines_13_ways_1_selComb;
    lines_14_ways_0_sel <= lines_14_ways_0_selComb;
    lines_14_ways_1_sel <= lines_14_ways_1_selComb;
    lines_15_ways_0_sel <= lines_15_ways_0_selComb;
    lines_15_ways_1_sel <= lines_15_ways_1_selComb;
    if(compaction_moveIt) begin
      lines_0_ways_0_context_staticWake <= lines_1_ways_0_context_staticWake;
      lines_0_ways_0_context_physRd <= lines_1_ways_0_context_physRd;
      lines_0_ways_0_context_robId <= lines_1_ways_0_context_robId;
      lines_0_ways_0_context_euCtx_0 <= lines_1_ways_0_context_euCtx_0;
      lines_0_ways_0_context_euCtx_1 <= lines_1_ways_0_context_euCtx_1;
      lines_0_ways_0_triggers <= (lines_1_ways_0_triggers >>> 2'd2);
      lines_0_ways_0_sel <= lines_1_ways_0_selComb;
      lines_0_ways_1_context_staticWake <= lines_1_ways_1_context_staticWake;
      lines_0_ways_1_context_physRd <= lines_1_ways_1_context_physRd;
      lines_0_ways_1_context_robId <= lines_1_ways_1_context_robId;
      lines_0_ways_1_context_euCtx_0 <= lines_1_ways_1_context_euCtx_0;
      lines_0_ways_1_context_euCtx_1 <= lines_1_ways_1_context_euCtx_1;
      lines_0_ways_1_triggers <= (lines_1_ways_1_triggers >>> 2'd2);
      lines_0_ways_1_sel <= lines_1_ways_1_selComb;
      lines_1_ways_0_context_staticWake <= lines_2_ways_0_context_staticWake;
      lines_1_ways_0_context_physRd <= lines_2_ways_0_context_physRd;
      lines_1_ways_0_context_robId <= lines_2_ways_0_context_robId;
      lines_1_ways_0_context_euCtx_0 <= lines_2_ways_0_context_euCtx_0;
      lines_1_ways_0_context_euCtx_1 <= lines_2_ways_0_context_euCtx_1;
      lines_1_ways_0_triggers <= (lines_2_ways_0_triggers >>> 2'd2);
      lines_1_ways_0_sel <= lines_2_ways_0_selComb;
      lines_1_ways_1_context_staticWake <= lines_2_ways_1_context_staticWake;
      lines_1_ways_1_context_physRd <= lines_2_ways_1_context_physRd;
      lines_1_ways_1_context_robId <= lines_2_ways_1_context_robId;
      lines_1_ways_1_context_euCtx_0 <= lines_2_ways_1_context_euCtx_0;
      lines_1_ways_1_context_euCtx_1 <= lines_2_ways_1_context_euCtx_1;
      lines_1_ways_1_triggers <= (lines_2_ways_1_triggers >>> 2'd2);
      lines_1_ways_1_sel <= lines_2_ways_1_selComb;
      lines_2_ways_0_context_staticWake <= lines_3_ways_0_context_staticWake;
      lines_2_ways_0_context_physRd <= lines_3_ways_0_context_physRd;
      lines_2_ways_0_context_robId <= lines_3_ways_0_context_robId;
      lines_2_ways_0_context_euCtx_0 <= lines_3_ways_0_context_euCtx_0;
      lines_2_ways_0_context_euCtx_1 <= lines_3_ways_0_context_euCtx_1;
      lines_2_ways_0_triggers <= (lines_3_ways_0_triggers >>> 2'd2);
      lines_2_ways_0_sel <= lines_3_ways_0_selComb;
      lines_2_ways_1_context_staticWake <= lines_3_ways_1_context_staticWake;
      lines_2_ways_1_context_physRd <= lines_3_ways_1_context_physRd;
      lines_2_ways_1_context_robId <= lines_3_ways_1_context_robId;
      lines_2_ways_1_context_euCtx_0 <= lines_3_ways_1_context_euCtx_0;
      lines_2_ways_1_context_euCtx_1 <= lines_3_ways_1_context_euCtx_1;
      lines_2_ways_1_triggers <= (lines_3_ways_1_triggers >>> 2'd2);
      lines_2_ways_1_sel <= lines_3_ways_1_selComb;
      lines_3_ways_0_context_staticWake <= lines_4_ways_0_context_staticWake;
      lines_3_ways_0_context_physRd <= lines_4_ways_0_context_physRd;
      lines_3_ways_0_context_robId <= lines_4_ways_0_context_robId;
      lines_3_ways_0_context_euCtx_0 <= lines_4_ways_0_context_euCtx_0;
      lines_3_ways_0_context_euCtx_1 <= lines_4_ways_0_context_euCtx_1;
      lines_3_ways_0_triggers <= (lines_4_ways_0_triggers >>> 2'd2);
      lines_3_ways_0_sel <= lines_4_ways_0_selComb;
      lines_3_ways_1_context_staticWake <= lines_4_ways_1_context_staticWake;
      lines_3_ways_1_context_physRd <= lines_4_ways_1_context_physRd;
      lines_3_ways_1_context_robId <= lines_4_ways_1_context_robId;
      lines_3_ways_1_context_euCtx_0 <= lines_4_ways_1_context_euCtx_0;
      lines_3_ways_1_context_euCtx_1 <= lines_4_ways_1_context_euCtx_1;
      lines_3_ways_1_triggers <= (lines_4_ways_1_triggers >>> 2'd2);
      lines_3_ways_1_sel <= lines_4_ways_1_selComb;
      lines_4_ways_0_context_staticWake <= lines_5_ways_0_context_staticWake;
      lines_4_ways_0_context_physRd <= lines_5_ways_0_context_physRd;
      lines_4_ways_0_context_robId <= lines_5_ways_0_context_robId;
      lines_4_ways_0_context_euCtx_0 <= lines_5_ways_0_context_euCtx_0;
      lines_4_ways_0_context_euCtx_1 <= lines_5_ways_0_context_euCtx_1;
      lines_4_ways_0_triggers <= (lines_5_ways_0_triggers >>> 2'd2);
      lines_4_ways_0_sel <= lines_5_ways_0_selComb;
      lines_4_ways_1_context_staticWake <= lines_5_ways_1_context_staticWake;
      lines_4_ways_1_context_physRd <= lines_5_ways_1_context_physRd;
      lines_4_ways_1_context_robId <= lines_5_ways_1_context_robId;
      lines_4_ways_1_context_euCtx_0 <= lines_5_ways_1_context_euCtx_0;
      lines_4_ways_1_context_euCtx_1 <= lines_5_ways_1_context_euCtx_1;
      lines_4_ways_1_triggers <= (lines_5_ways_1_triggers >>> 2'd2);
      lines_4_ways_1_sel <= lines_5_ways_1_selComb;
      lines_5_ways_0_context_staticWake <= lines_6_ways_0_context_staticWake;
      lines_5_ways_0_context_physRd <= lines_6_ways_0_context_physRd;
      lines_5_ways_0_context_robId <= lines_6_ways_0_context_robId;
      lines_5_ways_0_context_euCtx_0 <= lines_6_ways_0_context_euCtx_0;
      lines_5_ways_0_context_euCtx_1 <= lines_6_ways_0_context_euCtx_1;
      lines_5_ways_0_triggers <= (lines_6_ways_0_triggers >>> 2'd2);
      lines_5_ways_0_sel <= lines_6_ways_0_selComb;
      lines_5_ways_1_context_staticWake <= lines_6_ways_1_context_staticWake;
      lines_5_ways_1_context_physRd <= lines_6_ways_1_context_physRd;
      lines_5_ways_1_context_robId <= lines_6_ways_1_context_robId;
      lines_5_ways_1_context_euCtx_0 <= lines_6_ways_1_context_euCtx_0;
      lines_5_ways_1_context_euCtx_1 <= lines_6_ways_1_context_euCtx_1;
      lines_5_ways_1_triggers <= (lines_6_ways_1_triggers >>> 2'd2);
      lines_5_ways_1_sel <= lines_6_ways_1_selComb;
      lines_6_ways_0_context_staticWake <= lines_7_ways_0_context_staticWake;
      lines_6_ways_0_context_physRd <= lines_7_ways_0_context_physRd;
      lines_6_ways_0_context_robId <= lines_7_ways_0_context_robId;
      lines_6_ways_0_context_euCtx_0 <= lines_7_ways_0_context_euCtx_0;
      lines_6_ways_0_context_euCtx_1 <= lines_7_ways_0_context_euCtx_1;
      lines_6_ways_0_triggers <= (lines_7_ways_0_triggers >>> 2'd2);
      lines_6_ways_0_sel <= lines_7_ways_0_selComb;
      lines_6_ways_1_context_staticWake <= lines_7_ways_1_context_staticWake;
      lines_6_ways_1_context_physRd <= lines_7_ways_1_context_physRd;
      lines_6_ways_1_context_robId <= lines_7_ways_1_context_robId;
      lines_6_ways_1_context_euCtx_0 <= lines_7_ways_1_context_euCtx_0;
      lines_6_ways_1_context_euCtx_1 <= lines_7_ways_1_context_euCtx_1;
      lines_6_ways_1_triggers <= (lines_7_ways_1_triggers >>> 2'd2);
      lines_6_ways_1_sel <= lines_7_ways_1_selComb;
      lines_7_ways_0_context_staticWake <= lines_8_ways_0_context_staticWake;
      lines_7_ways_0_context_physRd <= lines_8_ways_0_context_physRd;
      lines_7_ways_0_context_robId <= lines_8_ways_0_context_robId;
      lines_7_ways_0_context_euCtx_0 <= lines_8_ways_0_context_euCtx_0;
      lines_7_ways_0_context_euCtx_1 <= lines_8_ways_0_context_euCtx_1;
      lines_7_ways_0_triggers <= (lines_8_ways_0_triggers >>> 2'd2);
      lines_7_ways_0_sel <= lines_8_ways_0_selComb;
      lines_7_ways_1_context_staticWake <= lines_8_ways_1_context_staticWake;
      lines_7_ways_1_context_physRd <= lines_8_ways_1_context_physRd;
      lines_7_ways_1_context_robId <= lines_8_ways_1_context_robId;
      lines_7_ways_1_context_euCtx_0 <= lines_8_ways_1_context_euCtx_0;
      lines_7_ways_1_context_euCtx_1 <= lines_8_ways_1_context_euCtx_1;
      lines_7_ways_1_triggers <= (lines_8_ways_1_triggers >>> 2'd2);
      lines_7_ways_1_sel <= lines_8_ways_1_selComb;
      lines_8_ways_0_context_staticWake <= lines_9_ways_0_context_staticWake;
      lines_8_ways_0_context_physRd <= lines_9_ways_0_context_physRd;
      lines_8_ways_0_context_robId <= lines_9_ways_0_context_robId;
      lines_8_ways_0_context_euCtx_0 <= lines_9_ways_0_context_euCtx_0;
      lines_8_ways_0_context_euCtx_1 <= lines_9_ways_0_context_euCtx_1;
      lines_8_ways_0_triggers <= (lines_9_ways_0_triggers >>> 2'd2);
      lines_8_ways_0_sel <= lines_9_ways_0_selComb;
      lines_8_ways_1_context_staticWake <= lines_9_ways_1_context_staticWake;
      lines_8_ways_1_context_physRd <= lines_9_ways_1_context_physRd;
      lines_8_ways_1_context_robId <= lines_9_ways_1_context_robId;
      lines_8_ways_1_context_euCtx_0 <= lines_9_ways_1_context_euCtx_0;
      lines_8_ways_1_context_euCtx_1 <= lines_9_ways_1_context_euCtx_1;
      lines_8_ways_1_triggers <= (lines_9_ways_1_triggers >>> 2'd2);
      lines_8_ways_1_sel <= lines_9_ways_1_selComb;
      lines_9_ways_0_context_staticWake <= lines_10_ways_0_context_staticWake;
      lines_9_ways_0_context_physRd <= lines_10_ways_0_context_physRd;
      lines_9_ways_0_context_robId <= lines_10_ways_0_context_robId;
      lines_9_ways_0_context_euCtx_0 <= lines_10_ways_0_context_euCtx_0;
      lines_9_ways_0_context_euCtx_1 <= lines_10_ways_0_context_euCtx_1;
      lines_9_ways_0_triggers <= (lines_10_ways_0_triggers >>> 2'd2);
      lines_9_ways_0_sel <= lines_10_ways_0_selComb;
      lines_9_ways_1_context_staticWake <= lines_10_ways_1_context_staticWake;
      lines_9_ways_1_context_physRd <= lines_10_ways_1_context_physRd;
      lines_9_ways_1_context_robId <= lines_10_ways_1_context_robId;
      lines_9_ways_1_context_euCtx_0 <= lines_10_ways_1_context_euCtx_0;
      lines_9_ways_1_context_euCtx_1 <= lines_10_ways_1_context_euCtx_1;
      lines_9_ways_1_triggers <= (lines_10_ways_1_triggers >>> 2'd2);
      lines_9_ways_1_sel <= lines_10_ways_1_selComb;
      lines_10_ways_0_context_staticWake <= lines_11_ways_0_context_staticWake;
      lines_10_ways_0_context_physRd <= lines_11_ways_0_context_physRd;
      lines_10_ways_0_context_robId <= lines_11_ways_0_context_robId;
      lines_10_ways_0_context_euCtx_0 <= lines_11_ways_0_context_euCtx_0;
      lines_10_ways_0_context_euCtx_1 <= lines_11_ways_0_context_euCtx_1;
      lines_10_ways_0_triggers <= (lines_11_ways_0_triggers >>> 2'd2);
      lines_10_ways_0_sel <= lines_11_ways_0_selComb;
      lines_10_ways_1_context_staticWake <= lines_11_ways_1_context_staticWake;
      lines_10_ways_1_context_physRd <= lines_11_ways_1_context_physRd;
      lines_10_ways_1_context_robId <= lines_11_ways_1_context_robId;
      lines_10_ways_1_context_euCtx_0 <= lines_11_ways_1_context_euCtx_0;
      lines_10_ways_1_context_euCtx_1 <= lines_11_ways_1_context_euCtx_1;
      lines_10_ways_1_triggers <= (lines_11_ways_1_triggers >>> 2'd2);
      lines_10_ways_1_sel <= lines_11_ways_1_selComb;
      lines_11_ways_0_context_staticWake <= lines_12_ways_0_context_staticWake;
      lines_11_ways_0_context_physRd <= lines_12_ways_0_context_physRd;
      lines_11_ways_0_context_robId <= lines_12_ways_0_context_robId;
      lines_11_ways_0_context_euCtx_0 <= lines_12_ways_0_context_euCtx_0;
      lines_11_ways_0_context_euCtx_1 <= lines_12_ways_0_context_euCtx_1;
      lines_11_ways_0_triggers <= (lines_12_ways_0_triggers >>> 2'd2);
      lines_11_ways_0_sel <= lines_12_ways_0_selComb;
      lines_11_ways_1_context_staticWake <= lines_12_ways_1_context_staticWake;
      lines_11_ways_1_context_physRd <= lines_12_ways_1_context_physRd;
      lines_11_ways_1_context_robId <= lines_12_ways_1_context_robId;
      lines_11_ways_1_context_euCtx_0 <= lines_12_ways_1_context_euCtx_0;
      lines_11_ways_1_context_euCtx_1 <= lines_12_ways_1_context_euCtx_1;
      lines_11_ways_1_triggers <= (lines_12_ways_1_triggers >>> 2'd2);
      lines_11_ways_1_sel <= lines_12_ways_1_selComb;
      lines_12_ways_0_context_staticWake <= lines_13_ways_0_context_staticWake;
      lines_12_ways_0_context_physRd <= lines_13_ways_0_context_physRd;
      lines_12_ways_0_context_robId <= lines_13_ways_0_context_robId;
      lines_12_ways_0_context_euCtx_0 <= lines_13_ways_0_context_euCtx_0;
      lines_12_ways_0_context_euCtx_1 <= lines_13_ways_0_context_euCtx_1;
      lines_12_ways_0_triggers <= (lines_13_ways_0_triggers >>> 2'd2);
      lines_12_ways_0_sel <= lines_13_ways_0_selComb;
      lines_12_ways_1_context_staticWake <= lines_13_ways_1_context_staticWake;
      lines_12_ways_1_context_physRd <= lines_13_ways_1_context_physRd;
      lines_12_ways_1_context_robId <= lines_13_ways_1_context_robId;
      lines_12_ways_1_context_euCtx_0 <= lines_13_ways_1_context_euCtx_0;
      lines_12_ways_1_context_euCtx_1 <= lines_13_ways_1_context_euCtx_1;
      lines_12_ways_1_triggers <= (lines_13_ways_1_triggers >>> 2'd2);
      lines_12_ways_1_sel <= lines_13_ways_1_selComb;
      lines_13_ways_0_context_staticWake <= lines_14_ways_0_context_staticWake;
      lines_13_ways_0_context_physRd <= lines_14_ways_0_context_physRd;
      lines_13_ways_0_context_robId <= lines_14_ways_0_context_robId;
      lines_13_ways_0_context_euCtx_0 <= lines_14_ways_0_context_euCtx_0;
      lines_13_ways_0_context_euCtx_1 <= lines_14_ways_0_context_euCtx_1;
      lines_13_ways_0_triggers <= (lines_14_ways_0_triggers >>> 2'd2);
      lines_13_ways_0_sel <= lines_14_ways_0_selComb;
      lines_13_ways_1_context_staticWake <= lines_14_ways_1_context_staticWake;
      lines_13_ways_1_context_physRd <= lines_14_ways_1_context_physRd;
      lines_13_ways_1_context_robId <= lines_14_ways_1_context_robId;
      lines_13_ways_1_context_euCtx_0 <= lines_14_ways_1_context_euCtx_0;
      lines_13_ways_1_context_euCtx_1 <= lines_14_ways_1_context_euCtx_1;
      lines_13_ways_1_triggers <= (lines_14_ways_1_triggers >>> 2'd2);
      lines_13_ways_1_sel <= lines_14_ways_1_selComb;
      lines_14_ways_0_context_staticWake <= lines_15_ways_0_context_staticWake;
      lines_14_ways_0_context_physRd <= lines_15_ways_0_context_physRd;
      lines_14_ways_0_context_robId <= lines_15_ways_0_context_robId;
      lines_14_ways_0_context_euCtx_0 <= lines_15_ways_0_context_euCtx_0;
      lines_14_ways_0_context_euCtx_1 <= lines_15_ways_0_context_euCtx_1;
      lines_14_ways_0_triggers <= (lines_15_ways_0_triggers >>> 2'd2);
      lines_14_ways_0_sel <= lines_15_ways_0_selComb;
      lines_14_ways_1_context_staticWake <= lines_15_ways_1_context_staticWake;
      lines_14_ways_1_context_physRd <= lines_15_ways_1_context_physRd;
      lines_14_ways_1_context_robId <= lines_15_ways_1_context_robId;
      lines_14_ways_1_context_euCtx_0 <= lines_15_ways_1_context_euCtx_0;
      lines_14_ways_1_context_euCtx_1 <= lines_15_ways_1_context_euCtx_1;
      lines_14_ways_1_triggers <= (lines_15_ways_1_triggers >>> 2'd2);
      lines_14_ways_1_sel <= lines_15_ways_1_selComb;
      lines_15_ways_0_context_staticWake <= io_push_payload_slots_0_context_staticWake;
      lines_15_ways_0_context_physRd <= io_push_payload_slots_0_context_physRd;
      lines_15_ways_0_context_robId <= io_push_payload_slots_0_context_robId;
      lines_15_ways_0_context_euCtx_0 <= io_push_payload_slots_0_context_euCtx_0;
      lines_15_ways_0_context_euCtx_1 <= io_push_payload_slots_0_context_euCtx_1;
      lines_15_ways_0_triggers <= io_push_payload_slots_0_event[30:0];
      lines_15_ways_0_sel <= io_push_payload_slots_0_sel;
      lines_15_ways_1_context_staticWake <= io_push_payload_slots_1_context_staticWake;
      lines_15_ways_1_context_physRd <= io_push_payload_slots_1_context_physRd;
      lines_15_ways_1_context_robId <= io_push_payload_slots_1_context_robId;
      lines_15_ways_1_context_euCtx_0 <= io_push_payload_slots_1_context_euCtx_0;
      lines_15_ways_1_context_euCtx_1 <= io_push_payload_slots_1_context_euCtx_1;
      lines_15_ways_1_triggers <= io_push_payload_slots_1_event;
      lines_15_ways_1_sel <= io_push_payload_slots_1_sel;
    end
    if(when_IssueQueue_l109) begin
      lines_0_ways_0_triggers[0] <= 1'b0;
      lines_0_ways_1_triggers[0] <= 1'b0;
      lines_1_ways_0_triggers[0] <= 1'b0;
      lines_1_ways_1_triggers[0] <= 1'b0;
      lines_2_ways_0_triggers[0] <= 1'b0;
      lines_2_ways_1_triggers[0] <= 1'b0;
      lines_3_ways_0_triggers[0] <= 1'b0;
      lines_3_ways_1_triggers[0] <= 1'b0;
      lines_4_ways_0_triggers[0] <= 1'b0;
      lines_4_ways_1_triggers[0] <= 1'b0;
      lines_5_ways_0_triggers[0] <= 1'b0;
      lines_5_ways_1_triggers[0] <= 1'b0;
      lines_6_ways_0_triggers[0] <= 1'b0;
      lines_6_ways_1_triggers[0] <= 1'b0;
      lines_7_ways_0_triggers[0] <= 1'b0;
      lines_7_ways_1_triggers[0] <= 1'b0;
      lines_8_ways_0_triggers[0] <= 1'b0;
      lines_8_ways_1_triggers[0] <= 1'b0;
      lines_9_ways_0_triggers[0] <= 1'b0;
      lines_9_ways_1_triggers[0] <= 1'b0;
      lines_10_ways_0_triggers[0] <= 1'b0;
      lines_10_ways_1_triggers[0] <= 1'b0;
      lines_11_ways_0_triggers[0] <= 1'b0;
      lines_11_ways_1_triggers[0] <= 1'b0;
      lines_12_ways_0_triggers[0] <= 1'b0;
      lines_12_ways_1_triggers[0] <= 1'b0;
      lines_13_ways_0_triggers[0] <= 1'b0;
      lines_13_ways_1_triggers[0] <= 1'b0;
      lines_14_ways_0_triggers[0] <= 1'b0;
      lines_14_ways_1_triggers[0] <= 1'b0;
      lines_15_ways_0_triggers[0] <= 1'b0;
      lines_15_ways_1_triggers[0] <= 1'b0;
    end
    if(when_IssueQueue_l109_1) begin
      lines_0_ways_1_triggers[1] <= 1'b0;
      lines_1_ways_0_triggers[1] <= 1'b0;
      lines_1_ways_1_triggers[1] <= 1'b0;
      lines_2_ways_0_triggers[1] <= 1'b0;
      lines_2_ways_1_triggers[1] <= 1'b0;
      lines_3_ways_0_triggers[1] <= 1'b0;
      lines_3_ways_1_triggers[1] <= 1'b0;
      lines_4_ways_0_triggers[1] <= 1'b0;
      lines_4_ways_1_triggers[1] <= 1'b0;
      lines_5_ways_0_triggers[1] <= 1'b0;
      lines_5_ways_1_triggers[1] <= 1'b0;
      lines_6_ways_0_triggers[1] <= 1'b0;
      lines_6_ways_1_triggers[1] <= 1'b0;
      lines_7_ways_0_triggers[1] <= 1'b0;
      lines_7_ways_1_triggers[1] <= 1'b0;
      lines_8_ways_0_triggers[1] <= 1'b0;
      lines_8_ways_1_triggers[1] <= 1'b0;
      lines_9_ways_0_triggers[1] <= 1'b0;
      lines_9_ways_1_triggers[1] <= 1'b0;
      lines_10_ways_0_triggers[1] <= 1'b0;
      lines_10_ways_1_triggers[1] <= 1'b0;
      lines_11_ways_0_triggers[1] <= 1'b0;
      lines_11_ways_1_triggers[1] <= 1'b0;
      lines_12_ways_0_triggers[1] <= 1'b0;
      lines_12_ways_1_triggers[1] <= 1'b0;
      lines_13_ways_0_triggers[1] <= 1'b0;
      lines_13_ways_1_triggers[1] <= 1'b0;
      lines_14_ways_0_triggers[1] <= 1'b0;
      lines_14_ways_1_triggers[1] <= 1'b0;
      lines_15_ways_0_triggers[1] <= 1'b0;
      lines_15_ways_1_triggers[1] <= 1'b0;
    end
    if(when_IssueQueue_l109_2) begin
      lines_1_ways_0_triggers[2] <= 1'b0;
      lines_1_ways_1_triggers[2] <= 1'b0;
      lines_2_ways_0_triggers[2] <= 1'b0;
      lines_2_ways_1_triggers[2] <= 1'b0;
      lines_3_ways_0_triggers[2] <= 1'b0;
      lines_3_ways_1_triggers[2] <= 1'b0;
      lines_4_ways_0_triggers[2] <= 1'b0;
      lines_4_ways_1_triggers[2] <= 1'b0;
      lines_5_ways_0_triggers[2] <= 1'b0;
      lines_5_ways_1_triggers[2] <= 1'b0;
      lines_6_ways_0_triggers[2] <= 1'b0;
      lines_6_ways_1_triggers[2] <= 1'b0;
      lines_7_ways_0_triggers[2] <= 1'b0;
      lines_7_ways_1_triggers[2] <= 1'b0;
      lines_8_ways_0_triggers[2] <= 1'b0;
      lines_8_ways_1_triggers[2] <= 1'b0;
      lines_9_ways_0_triggers[2] <= 1'b0;
      lines_9_ways_1_triggers[2] <= 1'b0;
      lines_10_ways_0_triggers[2] <= 1'b0;
      lines_10_ways_1_triggers[2] <= 1'b0;
      lines_11_ways_0_triggers[2] <= 1'b0;
      lines_11_ways_1_triggers[2] <= 1'b0;
      lines_12_ways_0_triggers[2] <= 1'b0;
      lines_12_ways_1_triggers[2] <= 1'b0;
      lines_13_ways_0_triggers[2] <= 1'b0;
      lines_13_ways_1_triggers[2] <= 1'b0;
      lines_14_ways_0_triggers[2] <= 1'b0;
      lines_14_ways_1_triggers[2] <= 1'b0;
      lines_15_ways_0_triggers[2] <= 1'b0;
      lines_15_ways_1_triggers[2] <= 1'b0;
    end
    if(when_IssueQueue_l109_3) begin
      lines_1_ways_1_triggers[3] <= 1'b0;
      lines_2_ways_0_triggers[3] <= 1'b0;
      lines_2_ways_1_triggers[3] <= 1'b0;
      lines_3_ways_0_triggers[3] <= 1'b0;
      lines_3_ways_1_triggers[3] <= 1'b0;
      lines_4_ways_0_triggers[3] <= 1'b0;
      lines_4_ways_1_triggers[3] <= 1'b0;
      lines_5_ways_0_triggers[3] <= 1'b0;
      lines_5_ways_1_triggers[3] <= 1'b0;
      lines_6_ways_0_triggers[3] <= 1'b0;
      lines_6_ways_1_triggers[3] <= 1'b0;
      lines_7_ways_0_triggers[3] <= 1'b0;
      lines_7_ways_1_triggers[3] <= 1'b0;
      lines_8_ways_0_triggers[3] <= 1'b0;
      lines_8_ways_1_triggers[3] <= 1'b0;
      lines_9_ways_0_triggers[3] <= 1'b0;
      lines_9_ways_1_triggers[3] <= 1'b0;
      lines_10_ways_0_triggers[3] <= 1'b0;
      lines_10_ways_1_triggers[3] <= 1'b0;
      lines_11_ways_0_triggers[3] <= 1'b0;
      lines_11_ways_1_triggers[3] <= 1'b0;
      lines_12_ways_0_triggers[3] <= 1'b0;
      lines_12_ways_1_triggers[3] <= 1'b0;
      lines_13_ways_0_triggers[3] <= 1'b0;
      lines_13_ways_1_triggers[3] <= 1'b0;
      lines_14_ways_0_triggers[3] <= 1'b0;
      lines_14_ways_1_triggers[3] <= 1'b0;
      lines_15_ways_0_triggers[3] <= 1'b0;
      lines_15_ways_1_triggers[3] <= 1'b0;
    end
    if(when_IssueQueue_l109_4) begin
      lines_2_ways_0_triggers[4] <= 1'b0;
      lines_2_ways_1_triggers[4] <= 1'b0;
      lines_3_ways_0_triggers[4] <= 1'b0;
      lines_3_ways_1_triggers[4] <= 1'b0;
      lines_4_ways_0_triggers[4] <= 1'b0;
      lines_4_ways_1_triggers[4] <= 1'b0;
      lines_5_ways_0_triggers[4] <= 1'b0;
      lines_5_ways_1_triggers[4] <= 1'b0;
      lines_6_ways_0_triggers[4] <= 1'b0;
      lines_6_ways_1_triggers[4] <= 1'b0;
      lines_7_ways_0_triggers[4] <= 1'b0;
      lines_7_ways_1_triggers[4] <= 1'b0;
      lines_8_ways_0_triggers[4] <= 1'b0;
      lines_8_ways_1_triggers[4] <= 1'b0;
      lines_9_ways_0_triggers[4] <= 1'b0;
      lines_9_ways_1_triggers[4] <= 1'b0;
      lines_10_ways_0_triggers[4] <= 1'b0;
      lines_10_ways_1_triggers[4] <= 1'b0;
      lines_11_ways_0_triggers[4] <= 1'b0;
      lines_11_ways_1_triggers[4] <= 1'b0;
      lines_12_ways_0_triggers[4] <= 1'b0;
      lines_12_ways_1_triggers[4] <= 1'b0;
      lines_13_ways_0_triggers[4] <= 1'b0;
      lines_13_ways_1_triggers[4] <= 1'b0;
      lines_14_ways_0_triggers[4] <= 1'b0;
      lines_14_ways_1_triggers[4] <= 1'b0;
      lines_15_ways_0_triggers[4] <= 1'b0;
      lines_15_ways_1_triggers[4] <= 1'b0;
    end
    if(when_IssueQueue_l109_5) begin
      lines_2_ways_1_triggers[5] <= 1'b0;
      lines_3_ways_0_triggers[5] <= 1'b0;
      lines_3_ways_1_triggers[5] <= 1'b0;
      lines_4_ways_0_triggers[5] <= 1'b0;
      lines_4_ways_1_triggers[5] <= 1'b0;
      lines_5_ways_0_triggers[5] <= 1'b0;
      lines_5_ways_1_triggers[5] <= 1'b0;
      lines_6_ways_0_triggers[5] <= 1'b0;
      lines_6_ways_1_triggers[5] <= 1'b0;
      lines_7_ways_0_triggers[5] <= 1'b0;
      lines_7_ways_1_triggers[5] <= 1'b0;
      lines_8_ways_0_triggers[5] <= 1'b0;
      lines_8_ways_1_triggers[5] <= 1'b0;
      lines_9_ways_0_triggers[5] <= 1'b0;
      lines_9_ways_1_triggers[5] <= 1'b0;
      lines_10_ways_0_triggers[5] <= 1'b0;
      lines_10_ways_1_triggers[5] <= 1'b0;
      lines_11_ways_0_triggers[5] <= 1'b0;
      lines_11_ways_1_triggers[5] <= 1'b0;
      lines_12_ways_0_triggers[5] <= 1'b0;
      lines_12_ways_1_triggers[5] <= 1'b0;
      lines_13_ways_0_triggers[5] <= 1'b0;
      lines_13_ways_1_triggers[5] <= 1'b0;
      lines_14_ways_0_triggers[5] <= 1'b0;
      lines_14_ways_1_triggers[5] <= 1'b0;
      lines_15_ways_0_triggers[5] <= 1'b0;
      lines_15_ways_1_triggers[5] <= 1'b0;
    end
    if(when_IssueQueue_l109_6) begin
      lines_3_ways_0_triggers[6] <= 1'b0;
      lines_3_ways_1_triggers[6] <= 1'b0;
      lines_4_ways_0_triggers[6] <= 1'b0;
      lines_4_ways_1_triggers[6] <= 1'b0;
      lines_5_ways_0_triggers[6] <= 1'b0;
      lines_5_ways_1_triggers[6] <= 1'b0;
      lines_6_ways_0_triggers[6] <= 1'b0;
      lines_6_ways_1_triggers[6] <= 1'b0;
      lines_7_ways_0_triggers[6] <= 1'b0;
      lines_7_ways_1_triggers[6] <= 1'b0;
      lines_8_ways_0_triggers[6] <= 1'b0;
      lines_8_ways_1_triggers[6] <= 1'b0;
      lines_9_ways_0_triggers[6] <= 1'b0;
      lines_9_ways_1_triggers[6] <= 1'b0;
      lines_10_ways_0_triggers[6] <= 1'b0;
      lines_10_ways_1_triggers[6] <= 1'b0;
      lines_11_ways_0_triggers[6] <= 1'b0;
      lines_11_ways_1_triggers[6] <= 1'b0;
      lines_12_ways_0_triggers[6] <= 1'b0;
      lines_12_ways_1_triggers[6] <= 1'b0;
      lines_13_ways_0_triggers[6] <= 1'b0;
      lines_13_ways_1_triggers[6] <= 1'b0;
      lines_14_ways_0_triggers[6] <= 1'b0;
      lines_14_ways_1_triggers[6] <= 1'b0;
      lines_15_ways_0_triggers[6] <= 1'b0;
      lines_15_ways_1_triggers[6] <= 1'b0;
    end
    if(when_IssueQueue_l109_7) begin
      lines_3_ways_1_triggers[7] <= 1'b0;
      lines_4_ways_0_triggers[7] <= 1'b0;
      lines_4_ways_1_triggers[7] <= 1'b0;
      lines_5_ways_0_triggers[7] <= 1'b0;
      lines_5_ways_1_triggers[7] <= 1'b0;
      lines_6_ways_0_triggers[7] <= 1'b0;
      lines_6_ways_1_triggers[7] <= 1'b0;
      lines_7_ways_0_triggers[7] <= 1'b0;
      lines_7_ways_1_triggers[7] <= 1'b0;
      lines_8_ways_0_triggers[7] <= 1'b0;
      lines_8_ways_1_triggers[7] <= 1'b0;
      lines_9_ways_0_triggers[7] <= 1'b0;
      lines_9_ways_1_triggers[7] <= 1'b0;
      lines_10_ways_0_triggers[7] <= 1'b0;
      lines_10_ways_1_triggers[7] <= 1'b0;
      lines_11_ways_0_triggers[7] <= 1'b0;
      lines_11_ways_1_triggers[7] <= 1'b0;
      lines_12_ways_0_triggers[7] <= 1'b0;
      lines_12_ways_1_triggers[7] <= 1'b0;
      lines_13_ways_0_triggers[7] <= 1'b0;
      lines_13_ways_1_triggers[7] <= 1'b0;
      lines_14_ways_0_triggers[7] <= 1'b0;
      lines_14_ways_1_triggers[7] <= 1'b0;
      lines_15_ways_0_triggers[7] <= 1'b0;
      lines_15_ways_1_triggers[7] <= 1'b0;
    end
    if(when_IssueQueue_l109_8) begin
      lines_4_ways_0_triggers[8] <= 1'b0;
      lines_4_ways_1_triggers[8] <= 1'b0;
      lines_5_ways_0_triggers[8] <= 1'b0;
      lines_5_ways_1_triggers[8] <= 1'b0;
      lines_6_ways_0_triggers[8] <= 1'b0;
      lines_6_ways_1_triggers[8] <= 1'b0;
      lines_7_ways_0_triggers[8] <= 1'b0;
      lines_7_ways_1_triggers[8] <= 1'b0;
      lines_8_ways_0_triggers[8] <= 1'b0;
      lines_8_ways_1_triggers[8] <= 1'b0;
      lines_9_ways_0_triggers[8] <= 1'b0;
      lines_9_ways_1_triggers[8] <= 1'b0;
      lines_10_ways_0_triggers[8] <= 1'b0;
      lines_10_ways_1_triggers[8] <= 1'b0;
      lines_11_ways_0_triggers[8] <= 1'b0;
      lines_11_ways_1_triggers[8] <= 1'b0;
      lines_12_ways_0_triggers[8] <= 1'b0;
      lines_12_ways_1_triggers[8] <= 1'b0;
      lines_13_ways_0_triggers[8] <= 1'b0;
      lines_13_ways_1_triggers[8] <= 1'b0;
      lines_14_ways_0_triggers[8] <= 1'b0;
      lines_14_ways_1_triggers[8] <= 1'b0;
      lines_15_ways_0_triggers[8] <= 1'b0;
      lines_15_ways_1_triggers[8] <= 1'b0;
    end
    if(when_IssueQueue_l109_9) begin
      lines_4_ways_1_triggers[9] <= 1'b0;
      lines_5_ways_0_triggers[9] <= 1'b0;
      lines_5_ways_1_triggers[9] <= 1'b0;
      lines_6_ways_0_triggers[9] <= 1'b0;
      lines_6_ways_1_triggers[9] <= 1'b0;
      lines_7_ways_0_triggers[9] <= 1'b0;
      lines_7_ways_1_triggers[9] <= 1'b0;
      lines_8_ways_0_triggers[9] <= 1'b0;
      lines_8_ways_1_triggers[9] <= 1'b0;
      lines_9_ways_0_triggers[9] <= 1'b0;
      lines_9_ways_1_triggers[9] <= 1'b0;
      lines_10_ways_0_triggers[9] <= 1'b0;
      lines_10_ways_1_triggers[9] <= 1'b0;
      lines_11_ways_0_triggers[9] <= 1'b0;
      lines_11_ways_1_triggers[9] <= 1'b0;
      lines_12_ways_0_triggers[9] <= 1'b0;
      lines_12_ways_1_triggers[9] <= 1'b0;
      lines_13_ways_0_triggers[9] <= 1'b0;
      lines_13_ways_1_triggers[9] <= 1'b0;
      lines_14_ways_0_triggers[9] <= 1'b0;
      lines_14_ways_1_triggers[9] <= 1'b0;
      lines_15_ways_0_triggers[9] <= 1'b0;
      lines_15_ways_1_triggers[9] <= 1'b0;
    end
    if(when_IssueQueue_l109_10) begin
      lines_5_ways_0_triggers[10] <= 1'b0;
      lines_5_ways_1_triggers[10] <= 1'b0;
      lines_6_ways_0_triggers[10] <= 1'b0;
      lines_6_ways_1_triggers[10] <= 1'b0;
      lines_7_ways_0_triggers[10] <= 1'b0;
      lines_7_ways_1_triggers[10] <= 1'b0;
      lines_8_ways_0_triggers[10] <= 1'b0;
      lines_8_ways_1_triggers[10] <= 1'b0;
      lines_9_ways_0_triggers[10] <= 1'b0;
      lines_9_ways_1_triggers[10] <= 1'b0;
      lines_10_ways_0_triggers[10] <= 1'b0;
      lines_10_ways_1_triggers[10] <= 1'b0;
      lines_11_ways_0_triggers[10] <= 1'b0;
      lines_11_ways_1_triggers[10] <= 1'b0;
      lines_12_ways_0_triggers[10] <= 1'b0;
      lines_12_ways_1_triggers[10] <= 1'b0;
      lines_13_ways_0_triggers[10] <= 1'b0;
      lines_13_ways_1_triggers[10] <= 1'b0;
      lines_14_ways_0_triggers[10] <= 1'b0;
      lines_14_ways_1_triggers[10] <= 1'b0;
      lines_15_ways_0_triggers[10] <= 1'b0;
      lines_15_ways_1_triggers[10] <= 1'b0;
    end
    if(when_IssueQueue_l109_11) begin
      lines_5_ways_1_triggers[11] <= 1'b0;
      lines_6_ways_0_triggers[11] <= 1'b0;
      lines_6_ways_1_triggers[11] <= 1'b0;
      lines_7_ways_0_triggers[11] <= 1'b0;
      lines_7_ways_1_triggers[11] <= 1'b0;
      lines_8_ways_0_triggers[11] <= 1'b0;
      lines_8_ways_1_triggers[11] <= 1'b0;
      lines_9_ways_0_triggers[11] <= 1'b0;
      lines_9_ways_1_triggers[11] <= 1'b0;
      lines_10_ways_0_triggers[11] <= 1'b0;
      lines_10_ways_1_triggers[11] <= 1'b0;
      lines_11_ways_0_triggers[11] <= 1'b0;
      lines_11_ways_1_triggers[11] <= 1'b0;
      lines_12_ways_0_triggers[11] <= 1'b0;
      lines_12_ways_1_triggers[11] <= 1'b0;
      lines_13_ways_0_triggers[11] <= 1'b0;
      lines_13_ways_1_triggers[11] <= 1'b0;
      lines_14_ways_0_triggers[11] <= 1'b0;
      lines_14_ways_1_triggers[11] <= 1'b0;
      lines_15_ways_0_triggers[11] <= 1'b0;
      lines_15_ways_1_triggers[11] <= 1'b0;
    end
    if(when_IssueQueue_l109_12) begin
      lines_6_ways_0_triggers[12] <= 1'b0;
      lines_6_ways_1_triggers[12] <= 1'b0;
      lines_7_ways_0_triggers[12] <= 1'b0;
      lines_7_ways_1_triggers[12] <= 1'b0;
      lines_8_ways_0_triggers[12] <= 1'b0;
      lines_8_ways_1_triggers[12] <= 1'b0;
      lines_9_ways_0_triggers[12] <= 1'b0;
      lines_9_ways_1_triggers[12] <= 1'b0;
      lines_10_ways_0_triggers[12] <= 1'b0;
      lines_10_ways_1_triggers[12] <= 1'b0;
      lines_11_ways_0_triggers[12] <= 1'b0;
      lines_11_ways_1_triggers[12] <= 1'b0;
      lines_12_ways_0_triggers[12] <= 1'b0;
      lines_12_ways_1_triggers[12] <= 1'b0;
      lines_13_ways_0_triggers[12] <= 1'b0;
      lines_13_ways_1_triggers[12] <= 1'b0;
      lines_14_ways_0_triggers[12] <= 1'b0;
      lines_14_ways_1_triggers[12] <= 1'b0;
      lines_15_ways_0_triggers[12] <= 1'b0;
      lines_15_ways_1_triggers[12] <= 1'b0;
    end
    if(when_IssueQueue_l109_13) begin
      lines_6_ways_1_triggers[13] <= 1'b0;
      lines_7_ways_0_triggers[13] <= 1'b0;
      lines_7_ways_1_triggers[13] <= 1'b0;
      lines_8_ways_0_triggers[13] <= 1'b0;
      lines_8_ways_1_triggers[13] <= 1'b0;
      lines_9_ways_0_triggers[13] <= 1'b0;
      lines_9_ways_1_triggers[13] <= 1'b0;
      lines_10_ways_0_triggers[13] <= 1'b0;
      lines_10_ways_1_triggers[13] <= 1'b0;
      lines_11_ways_0_triggers[13] <= 1'b0;
      lines_11_ways_1_triggers[13] <= 1'b0;
      lines_12_ways_0_triggers[13] <= 1'b0;
      lines_12_ways_1_triggers[13] <= 1'b0;
      lines_13_ways_0_triggers[13] <= 1'b0;
      lines_13_ways_1_triggers[13] <= 1'b0;
      lines_14_ways_0_triggers[13] <= 1'b0;
      lines_14_ways_1_triggers[13] <= 1'b0;
      lines_15_ways_0_triggers[13] <= 1'b0;
      lines_15_ways_1_triggers[13] <= 1'b0;
    end
    if(when_IssueQueue_l109_14) begin
      lines_7_ways_0_triggers[14] <= 1'b0;
      lines_7_ways_1_triggers[14] <= 1'b0;
      lines_8_ways_0_triggers[14] <= 1'b0;
      lines_8_ways_1_triggers[14] <= 1'b0;
      lines_9_ways_0_triggers[14] <= 1'b0;
      lines_9_ways_1_triggers[14] <= 1'b0;
      lines_10_ways_0_triggers[14] <= 1'b0;
      lines_10_ways_1_triggers[14] <= 1'b0;
      lines_11_ways_0_triggers[14] <= 1'b0;
      lines_11_ways_1_triggers[14] <= 1'b0;
      lines_12_ways_0_triggers[14] <= 1'b0;
      lines_12_ways_1_triggers[14] <= 1'b0;
      lines_13_ways_0_triggers[14] <= 1'b0;
      lines_13_ways_1_triggers[14] <= 1'b0;
      lines_14_ways_0_triggers[14] <= 1'b0;
      lines_14_ways_1_triggers[14] <= 1'b0;
      lines_15_ways_0_triggers[14] <= 1'b0;
      lines_15_ways_1_triggers[14] <= 1'b0;
    end
    if(when_IssueQueue_l109_15) begin
      lines_7_ways_1_triggers[15] <= 1'b0;
      lines_8_ways_0_triggers[15] <= 1'b0;
      lines_8_ways_1_triggers[15] <= 1'b0;
      lines_9_ways_0_triggers[15] <= 1'b0;
      lines_9_ways_1_triggers[15] <= 1'b0;
      lines_10_ways_0_triggers[15] <= 1'b0;
      lines_10_ways_1_triggers[15] <= 1'b0;
      lines_11_ways_0_triggers[15] <= 1'b0;
      lines_11_ways_1_triggers[15] <= 1'b0;
      lines_12_ways_0_triggers[15] <= 1'b0;
      lines_12_ways_1_triggers[15] <= 1'b0;
      lines_13_ways_0_triggers[15] <= 1'b0;
      lines_13_ways_1_triggers[15] <= 1'b0;
      lines_14_ways_0_triggers[15] <= 1'b0;
      lines_14_ways_1_triggers[15] <= 1'b0;
      lines_15_ways_0_triggers[15] <= 1'b0;
      lines_15_ways_1_triggers[15] <= 1'b0;
    end
    if(when_IssueQueue_l109_16) begin
      lines_8_ways_0_triggers[16] <= 1'b0;
      lines_8_ways_1_triggers[16] <= 1'b0;
      lines_9_ways_0_triggers[16] <= 1'b0;
      lines_9_ways_1_triggers[16] <= 1'b0;
      lines_10_ways_0_triggers[16] <= 1'b0;
      lines_10_ways_1_triggers[16] <= 1'b0;
      lines_11_ways_0_triggers[16] <= 1'b0;
      lines_11_ways_1_triggers[16] <= 1'b0;
      lines_12_ways_0_triggers[16] <= 1'b0;
      lines_12_ways_1_triggers[16] <= 1'b0;
      lines_13_ways_0_triggers[16] <= 1'b0;
      lines_13_ways_1_triggers[16] <= 1'b0;
      lines_14_ways_0_triggers[16] <= 1'b0;
      lines_14_ways_1_triggers[16] <= 1'b0;
      lines_15_ways_0_triggers[16] <= 1'b0;
      lines_15_ways_1_triggers[16] <= 1'b0;
    end
    if(when_IssueQueue_l109_17) begin
      lines_8_ways_1_triggers[17] <= 1'b0;
      lines_9_ways_0_triggers[17] <= 1'b0;
      lines_9_ways_1_triggers[17] <= 1'b0;
      lines_10_ways_0_triggers[17] <= 1'b0;
      lines_10_ways_1_triggers[17] <= 1'b0;
      lines_11_ways_0_triggers[17] <= 1'b0;
      lines_11_ways_1_triggers[17] <= 1'b0;
      lines_12_ways_0_triggers[17] <= 1'b0;
      lines_12_ways_1_triggers[17] <= 1'b0;
      lines_13_ways_0_triggers[17] <= 1'b0;
      lines_13_ways_1_triggers[17] <= 1'b0;
      lines_14_ways_0_triggers[17] <= 1'b0;
      lines_14_ways_1_triggers[17] <= 1'b0;
      lines_15_ways_0_triggers[17] <= 1'b0;
      lines_15_ways_1_triggers[17] <= 1'b0;
    end
    if(when_IssueQueue_l109_18) begin
      lines_9_ways_0_triggers[18] <= 1'b0;
      lines_9_ways_1_triggers[18] <= 1'b0;
      lines_10_ways_0_triggers[18] <= 1'b0;
      lines_10_ways_1_triggers[18] <= 1'b0;
      lines_11_ways_0_triggers[18] <= 1'b0;
      lines_11_ways_1_triggers[18] <= 1'b0;
      lines_12_ways_0_triggers[18] <= 1'b0;
      lines_12_ways_1_triggers[18] <= 1'b0;
      lines_13_ways_0_triggers[18] <= 1'b0;
      lines_13_ways_1_triggers[18] <= 1'b0;
      lines_14_ways_0_triggers[18] <= 1'b0;
      lines_14_ways_1_triggers[18] <= 1'b0;
      lines_15_ways_0_triggers[18] <= 1'b0;
      lines_15_ways_1_triggers[18] <= 1'b0;
    end
    if(when_IssueQueue_l109_19) begin
      lines_9_ways_1_triggers[19] <= 1'b0;
      lines_10_ways_0_triggers[19] <= 1'b0;
      lines_10_ways_1_triggers[19] <= 1'b0;
      lines_11_ways_0_triggers[19] <= 1'b0;
      lines_11_ways_1_triggers[19] <= 1'b0;
      lines_12_ways_0_triggers[19] <= 1'b0;
      lines_12_ways_1_triggers[19] <= 1'b0;
      lines_13_ways_0_triggers[19] <= 1'b0;
      lines_13_ways_1_triggers[19] <= 1'b0;
      lines_14_ways_0_triggers[19] <= 1'b0;
      lines_14_ways_1_triggers[19] <= 1'b0;
      lines_15_ways_0_triggers[19] <= 1'b0;
      lines_15_ways_1_triggers[19] <= 1'b0;
    end
    if(when_IssueQueue_l109_20) begin
      lines_10_ways_0_triggers[20] <= 1'b0;
      lines_10_ways_1_triggers[20] <= 1'b0;
      lines_11_ways_0_triggers[20] <= 1'b0;
      lines_11_ways_1_triggers[20] <= 1'b0;
      lines_12_ways_0_triggers[20] <= 1'b0;
      lines_12_ways_1_triggers[20] <= 1'b0;
      lines_13_ways_0_triggers[20] <= 1'b0;
      lines_13_ways_1_triggers[20] <= 1'b0;
      lines_14_ways_0_triggers[20] <= 1'b0;
      lines_14_ways_1_triggers[20] <= 1'b0;
      lines_15_ways_0_triggers[20] <= 1'b0;
      lines_15_ways_1_triggers[20] <= 1'b0;
    end
    if(when_IssueQueue_l109_21) begin
      lines_10_ways_1_triggers[21] <= 1'b0;
      lines_11_ways_0_triggers[21] <= 1'b0;
      lines_11_ways_1_triggers[21] <= 1'b0;
      lines_12_ways_0_triggers[21] <= 1'b0;
      lines_12_ways_1_triggers[21] <= 1'b0;
      lines_13_ways_0_triggers[21] <= 1'b0;
      lines_13_ways_1_triggers[21] <= 1'b0;
      lines_14_ways_0_triggers[21] <= 1'b0;
      lines_14_ways_1_triggers[21] <= 1'b0;
      lines_15_ways_0_triggers[21] <= 1'b0;
      lines_15_ways_1_triggers[21] <= 1'b0;
    end
    if(when_IssueQueue_l109_22) begin
      lines_11_ways_0_triggers[22] <= 1'b0;
      lines_11_ways_1_triggers[22] <= 1'b0;
      lines_12_ways_0_triggers[22] <= 1'b0;
      lines_12_ways_1_triggers[22] <= 1'b0;
      lines_13_ways_0_triggers[22] <= 1'b0;
      lines_13_ways_1_triggers[22] <= 1'b0;
      lines_14_ways_0_triggers[22] <= 1'b0;
      lines_14_ways_1_triggers[22] <= 1'b0;
      lines_15_ways_0_triggers[22] <= 1'b0;
      lines_15_ways_1_triggers[22] <= 1'b0;
    end
    if(when_IssueQueue_l109_23) begin
      lines_11_ways_1_triggers[23] <= 1'b0;
      lines_12_ways_0_triggers[23] <= 1'b0;
      lines_12_ways_1_triggers[23] <= 1'b0;
      lines_13_ways_0_triggers[23] <= 1'b0;
      lines_13_ways_1_triggers[23] <= 1'b0;
      lines_14_ways_0_triggers[23] <= 1'b0;
      lines_14_ways_1_triggers[23] <= 1'b0;
      lines_15_ways_0_triggers[23] <= 1'b0;
      lines_15_ways_1_triggers[23] <= 1'b0;
    end
    if(when_IssueQueue_l109_24) begin
      lines_12_ways_0_triggers[24] <= 1'b0;
      lines_12_ways_1_triggers[24] <= 1'b0;
      lines_13_ways_0_triggers[24] <= 1'b0;
      lines_13_ways_1_triggers[24] <= 1'b0;
      lines_14_ways_0_triggers[24] <= 1'b0;
      lines_14_ways_1_triggers[24] <= 1'b0;
      lines_15_ways_0_triggers[24] <= 1'b0;
      lines_15_ways_1_triggers[24] <= 1'b0;
    end
    if(when_IssueQueue_l109_25) begin
      lines_12_ways_1_triggers[25] <= 1'b0;
      lines_13_ways_0_triggers[25] <= 1'b0;
      lines_13_ways_1_triggers[25] <= 1'b0;
      lines_14_ways_0_triggers[25] <= 1'b0;
      lines_14_ways_1_triggers[25] <= 1'b0;
      lines_15_ways_0_triggers[25] <= 1'b0;
      lines_15_ways_1_triggers[25] <= 1'b0;
    end
    if(when_IssueQueue_l109_26) begin
      lines_13_ways_0_triggers[26] <= 1'b0;
      lines_13_ways_1_triggers[26] <= 1'b0;
      lines_14_ways_0_triggers[26] <= 1'b0;
      lines_14_ways_1_triggers[26] <= 1'b0;
      lines_15_ways_0_triggers[26] <= 1'b0;
      lines_15_ways_1_triggers[26] <= 1'b0;
    end
    if(when_IssueQueue_l109_27) begin
      lines_13_ways_1_triggers[27] <= 1'b0;
      lines_14_ways_0_triggers[27] <= 1'b0;
      lines_14_ways_1_triggers[27] <= 1'b0;
      lines_15_ways_0_triggers[27] <= 1'b0;
      lines_15_ways_1_triggers[27] <= 1'b0;
    end
    if(when_IssueQueue_l109_28) begin
      lines_14_ways_0_triggers[28] <= 1'b0;
      lines_14_ways_1_triggers[28] <= 1'b0;
      lines_15_ways_0_triggers[28] <= 1'b0;
      lines_15_ways_1_triggers[28] <= 1'b0;
    end
    if(when_IssueQueue_l109_29) begin
      lines_14_ways_1_triggers[29] <= 1'b0;
      lines_15_ways_0_triggers[29] <= 1'b0;
      lines_15_ways_1_triggers[29] <= 1'b0;
    end
    if(when_IssueQueue_l109_30) begin
      lines_15_ways_0_triggers[30] <= 1'b0;
      lines_15_ways_1_triggers[30] <= 1'b0;
    end
    if(when_IssueQueue_l109_31) begin
      lines_15_ways_1_triggers[31] <= 1'b0;
    end
    if(clear) begin
      lines_0_ways_0_sel <= 2'b00;
      lines_0_ways_1_sel <= 2'b00;
      lines_1_ways_0_sel <= 2'b00;
      lines_1_ways_1_sel <= 2'b00;
      lines_2_ways_0_sel <= 2'b00;
      lines_2_ways_1_sel <= 2'b00;
      lines_3_ways_0_sel <= 2'b00;
      lines_3_ways_1_sel <= 2'b00;
      lines_4_ways_0_sel <= 2'b00;
      lines_4_ways_1_sel <= 2'b00;
      lines_5_ways_0_sel <= 2'b00;
      lines_5_ways_1_sel <= 2'b00;
      lines_6_ways_0_sel <= 2'b00;
      lines_6_ways_1_sel <= 2'b00;
      lines_7_ways_0_sel <= 2'b00;
      lines_7_ways_1_sel <= 2'b00;
      lines_8_ways_0_sel <= 2'b00;
      lines_8_ways_1_sel <= 2'b00;
      lines_9_ways_0_sel <= 2'b00;
      lines_9_ways_1_sel <= 2'b00;
      lines_10_ways_0_sel <= 2'b00;
      lines_10_ways_1_sel <= 2'b00;
      lines_11_ways_0_sel <= 2'b00;
      lines_11_ways_1_sel <= 2'b00;
      lines_12_ways_0_sel <= 2'b00;
      lines_12_ways_1_sel <= 2'b00;
      lines_13_ways_0_sel <= 2'b00;
      lines_13_ways_1_sel <= 2'b00;
      lines_14_ways_0_sel <= 2'b00;
      lines_14_ways_1_sel <= 2'b00;
      lines_15_ways_0_sel <= 2'b00;
      lines_15_ways_1_sel <= 2'b00;
    end
  end


endmodule

module PrefetchPredictor (
  input  wire          io_learn_valid,
  input  wire [31:0]   io_learn_payload_physical,
  input  wire          io_learn_payload_allocate,
  output wire          io_prediction_cmd_valid,
  input  wire          io_prediction_cmd_ready,
  output wire [31:0]   io_prediction_cmd_payload,
  input  wire          io_prediction_rsp_valid,
  input  wire          io_prediction_rsp_payload
);


  assign io_prediction_cmd_valid = 1'b0;
  assign io_prediction_cmd_payload = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;

endmodule

module DivRadix4 (
  input  wire          io_flush,
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [31:0]   io_cmd_payload_a,
  input  wire [31:0]   io_cmd_payload_b,
  output wire          io_rsp_valid,
  input  wire          io_rsp_ready,
  output wire [34:0]   io_rsp_payload_result,
  output wire [32:0]   io_rsp_payload_remain,
  input  wire          clk,
  input  wire          reset
);

  wire       [33:0]   _zz_div3;
  wire       [32:0]   _zz_div3_1;
  wire       [32:0]   _zz_div3_2;
  wire       [7:0]    _zz_shifter_1;
  wire       [15:0]   _zz_shifter_2;
  wire       [23:0]   _zz_shifter_3;
  reg        [3:0]    counter;
  reg                 busy;
  wire                io_rsp_fire;
  reg                 done;
  wire                when_DivRadix4_l32;
  reg        [31:0]   shifter;
  reg        [31:0]   numerator;
  reg        [31:0]   result;
  reg        [33:0]   div1;
  reg        [33:0]   div3;
  wire       [33:0]   div2;
  wire       [33:0]   shifted;
  wire       [34:0]   sub1;
  wire       [34:0]   sub2;
  wire       [34:0]   sub3;
  wire                when_DivRadix4_l51;
  reg        [33:0]   _zz_shifter;
  wire                when_DivRadix4_l55;
  wire                when_DivRadix4_l59;
  wire                when_DivRadix4_l63;
  wire                slicesZero_0;
  wire                slicesZero_1;
  wire                slicesZero_2;
  wire       [2:0]    shiftSel;
  wire       [3:0]    _zz_sel;
  wire                _zz_sel_1;
  wire                _zz_sel_2;
  wire                _zz_sel_3;
  reg        [3:0]    _zz_sel_4;
  wire       [3:0]    _zz_sel_5;
  wire                _zz_sel_6;
  wire                _zz_sel_7;
  wire                _zz_sel_8;
  wire       [1:0]    sel;
  wire                when_DivRadix4_l77;

  assign _zz_div3_1 = {1'b0,io_cmd_payload_b};
  assign _zz_div3 = {1'd0, _zz_div3_1};
  assign _zz_div3_2 = ({1'd0,io_cmd_payload_b} <<< 1'd1);
  assign _zz_shifter_1 = io_cmd_payload_a[31 : 24];
  assign _zz_shifter_2 = io_cmd_payload_a[31 : 16];
  assign _zz_shifter_3 = io_cmd_payload_a[31 : 8];
  assign io_rsp_fire = (io_rsp_valid && io_rsp_ready);
  assign when_DivRadix4_l32 = (busy && (counter == 4'b1111));
  assign div2 = (div1 <<< 1);
  assign shifted = {shifter,numerator[31 : 30]};
  assign sub1 = ({1'b0,shifted} - {1'b0,div1});
  assign sub2 = ({1'b0,shifted} - {1'b0,div2});
  assign sub3 = ({1'b0,shifted} - {1'b0,div3});
  assign io_rsp_valid = done;
  assign io_rsp_payload_result = {3'd0, result};
  assign io_rsp_payload_remain = {1'd0, shifter};
  assign io_cmd_ready = (! busy);
  assign when_DivRadix4_l51 = (! done);
  always @(*) begin
    _zz_shifter = shifted;
    if(when_DivRadix4_l55) begin
      _zz_shifter = sub1[33:0];
    end
    if(when_DivRadix4_l59) begin
      _zz_shifter = sub2[33:0];
    end
    if(when_DivRadix4_l63) begin
      _zz_shifter = sub3[33:0];
    end
  end

  assign when_DivRadix4_l55 = (! sub1[34]);
  assign when_DivRadix4_l59 = (! sub2[34]);
  assign when_DivRadix4_l63 = (! sub3[34]);
  assign slicesZero_0 = (io_cmd_payload_a[15 : 8] == 8'h00);
  assign slicesZero_1 = (io_cmd_payload_a[23 : 16] == 8'h00);
  assign slicesZero_2 = (io_cmd_payload_a[31 : 24] == 8'h00);
  assign shiftSel = {slicesZero_2,{(slicesZero_1 && slicesZero_2),((slicesZero_0 && slicesZero_1) && slicesZero_2)}};
  assign _zz_sel = {1'b1,shiftSel};
  assign _zz_sel_1 = _zz_sel[0];
  assign _zz_sel_2 = _zz_sel[1];
  assign _zz_sel_3 = _zz_sel[2];
  always @(*) begin
    _zz_sel_4[0] = (_zz_sel_1 && (! 1'b0));
    _zz_sel_4[1] = (_zz_sel_2 && (! _zz_sel_1));
    _zz_sel_4[2] = (_zz_sel_3 && (! ({_zz_sel_2,_zz_sel_1} != 2'b00)));
    _zz_sel_4[3] = (_zz_sel[3] && (! ({_zz_sel_3,{_zz_sel_2,_zz_sel_1}} != 3'b000)));
  end

  assign _zz_sel_5 = _zz_sel_4;
  assign _zz_sel_6 = _zz_sel_5[3];
  assign _zz_sel_7 = (_zz_sel_5[1] || _zz_sel_6);
  assign _zz_sel_8 = (_zz_sel_5[2] || _zz_sel_6);
  assign sel = {_zz_sel_8,_zz_sel_7};
  assign when_DivRadix4_l77 = (! busy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      busy <= 1'b0;
      done <= 1'b0;
    end else begin
      if(io_rsp_fire) begin
        busy <= 1'b0;
      end
      if(when_DivRadix4_l32) begin
        done <= 1'b1;
      end
      if(io_rsp_fire) begin
        done <= 1'b0;
      end
      if(when_DivRadix4_l77) begin
        busy <= io_cmd_valid;
      end
      if(io_flush) begin
        done <= 1'b0;
        busy <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(when_DivRadix4_l51) begin
      counter <= (counter + 4'b0001);
      result <= (result <<< 2);
      if(when_DivRadix4_l55) begin
        result[1 : 0] <= 2'b01;
      end
      if(when_DivRadix4_l59) begin
        result[1 : 0] <= 2'b10;
      end
      if(when_DivRadix4_l63) begin
        result[1 : 0] <= 2'b11;
      end
      shifter <= _zz_shifter[31:0];
      numerator <= (numerator <<< 2);
    end
    if(when_DivRadix4_l77) begin
      div1 <= {2'd0, io_cmd_payload_b};
      div3 <= (_zz_div3 + {1'b0,_zz_div3_2});
      result <= ((io_cmd_payload_b == 32'h00000000) ? 32'hffffffff : 32'h00000000);
      case(sel)
        2'b11 : begin
          counter <= 4'b0000;
          shifter <= 32'h00000000;
          numerator <= (io_cmd_payload_a <<< 0);
        end
        2'b10 : begin
          counter <= 4'b0100;
          shifter <= {24'd0, _zz_shifter_1};
          numerator <= (io_cmd_payload_a <<< 8);
        end
        2'b01 : begin
          counter <= 4'b1000;
          shifter <= {16'd0, _zz_shifter_2};
          numerator <= (io_cmd_payload_a <<< 16);
        end
        default : begin
          counter <= 4'b1100;
          shifter <= {8'd0, _zz_shifter_3};
          numerator <= (io_cmd_payload_a <<< 24);
        end
      endcase
    end
  end


endmodule

module StreamFifoLowLatency (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [5:0]    io_push_payload_robId,
  input  wire [1:0]    io_push_payload_mask,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [5:0]    io_pop_payload_robId,
  output wire [1:0]    io_pop_payload_mask,
  input  wire          io_flush,
  output wire [5:0]    io_occupancy,
  output wire [5:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  wire                fifo_io_push_ready;
  wire                fifo_io_pop_valid;
  wire       [5:0]    fifo_io_pop_payload_robId;
  wire       [1:0]    fifo_io_pop_payload_mask;
  wire       [5:0]    fifo_io_occupancy;
  wire       [5:0]    fifo_io_availability;

  StreamFifo fifo (
    .io_push_valid         (io_push_valid                 ), //i
    .io_push_ready         (fifo_io_push_ready            ), //o
    .io_push_payload_robId (io_push_payload_robId[5:0]    ), //i
    .io_push_payload_mask  (io_push_payload_mask[1:0]     ), //i
    .io_pop_valid          (fifo_io_pop_valid             ), //o
    .io_pop_ready          (io_pop_ready                  ), //i
    .io_pop_payload_robId  (fifo_io_pop_payload_robId[5:0]), //o
    .io_pop_payload_mask   (fifo_io_pop_payload_mask[1:0] ), //o
    .io_flush              (io_flush                      ), //i
    .io_occupancy          (fifo_io_occupancy[5:0]        ), //o
    .io_availability       (fifo_io_availability[5:0]     ), //o
    .clk                   (clk                           ), //i
    .reset                 (reset                         )  //i
  );
  assign io_push_ready = fifo_io_push_ready;
  assign io_pop_valid = fifo_io_pop_valid;
  assign io_pop_payload_robId = fifo_io_pop_payload_robId;
  assign io_pop_payload_mask = fifo_io_pop_payload_mask;
  assign io_occupancy = fifo_io_occupancy;
  assign io_availability = fifo_io_availability;

endmodule

module DataCache (
  input  wire          io_lock_valid,
  input  wire [31:0]   io_lock_address,
  input  wire          io_load_cmd_valid,
  output wire          io_load_cmd_ready,
  input  wire [31:0]   io_load_cmd_payload_virtual,
  input  wire [1:0]    io_load_cmd_payload_size,
  input  wire          io_load_cmd_payload_redoOnDataHazard,
  input  wire          io_load_cmd_payload_unlocked,
  input  wire          io_load_cmd_payload_unique,
  input  wire [31:0]   io_load_translated_physical,
  input  wire          io_load_translated_abord,
  input  wire [2:0]    io_load_cancels,
  output wire          io_load_rsp_valid,
  output wire [31:0]   io_load_rsp_payload_data,
  output wire          io_load_rsp_payload_fault,
  output wire          io_load_rsp_payload_redo,
  output wire [1:0]    io_load_rsp_payload_refillSlot,
  output wire          io_load_rsp_payload_refillSlotAny,
  input  wire          io_store_cmd_valid,
  output wire          io_store_cmd_ready,
  input  wire [31:0]   io_store_cmd_payload_address,
  input  wire [31:0]   io_store_cmd_payload_data,
  input  wire [3:0]    io_store_cmd_payload_mask,
  input  wire          io_store_cmd_payload_generation,
  input  wire          io_store_cmd_payload_io,
  input  wire          io_store_cmd_payload_flush,
  input  wire          io_store_cmd_payload_flushFree,
  input  wire          io_store_cmd_payload_prefetch,
  output wire          io_store_rsp_valid,
  output wire          io_store_rsp_payload_fault,
  output wire          io_store_rsp_payload_redo,
  output wire [1:0]    io_store_rsp_payload_refillSlot,
  output wire          io_store_rsp_payload_refillSlotAny,
  output wire          io_store_rsp_payload_generationKo,
  output wire          io_store_rsp_payload_flush,
  output wire          io_store_rsp_payload_prefetch,
  output wire [31:0]   io_store_rsp_payload_address,
  output wire          io_store_rsp_payload_io,
  output wire          io_mem_read_cmd_valid,
  input  wire          io_mem_read_cmd_ready,
  output wire [0:0]    io_mem_read_cmd_payload_id,
  output wire [31:0]   io_mem_read_cmd_payload_address,
  input  wire          io_mem_read_rsp_valid,
  output wire          io_mem_read_rsp_ready,
  input  wire [0:0]    io_mem_read_rsp_payload_id,
  input  wire [63:0]   io_mem_read_rsp_payload_data,
  input  wire          io_mem_read_rsp_payload_error,
  output wire          io_mem_write_cmd_valid,
  input  wire          io_mem_write_cmd_ready,
  output wire          io_mem_write_cmd_payload_last,
  output wire [31:0]   io_mem_write_cmd_payload_fragment_address,
  output wire [63:0]   io_mem_write_cmd_payload_fragment_data,
  output wire [0:0]    io_mem_write_cmd_payload_fragment_id,
  input  wire          io_mem_write_rsp_valid,
  input  wire          io_mem_write_rsp_payload_error,
  input  wire [0:0]    io_mem_write_rsp_payload_id,
  output reg  [1:0]    io_refillCompletions,
  output wire          io_refillEvent,
  output wire          io_writebackEvent,
  output wire          io_writebackBusy,
  output wire          io_tagEvent,
  input  wire          clk,
  input  wire          reset
);

  reg        [63:0]   _zz_banks_0_mem_port1;
  reg        [63:0]   _zz_banks_1_mem_port1;
  reg        [63:0]   _zz_banks_2_mem_port1;
  reg        [63:0]   _zz_banks_3_mem_port1;
  wire       [21:0]   _zz_ways_0_mem_port1;
  wire       [21:0]   _zz_ways_0_mem_port2;
  wire       [21:0]   _zz_ways_1_mem_port1;
  wire       [21:0]   _zz_ways_1_mem_port2;
  wire       [21:0]   _zz_ways_2_mem_port1;
  wire       [21:0]   _zz_ways_2_mem_port2;
  wire       [21:0]   _zz_ways_3_mem_port1;
  wire       [21:0]   _zz_ways_3_mem_port2;
  wire       [3:0]    _zz_status_mem_port1;
  wire       [3:0]    _zz_status_mem_port2;
  wire       [2:0]    _zz_plru_ram_port1;
  wire       [2:0]    _zz_plru_ram_port2;
  reg        [63:0]   _zz_writeback_victimBuffer_port1;
  wire       [21:0]   _zz_ways_0_mem_port;
  wire                _zz_ways_0_mem_port_1;
  wire       [21:0]   _zz_ways_1_mem_port;
  wire                _zz_ways_1_mem_port_1;
  wire       [21:0]   _zz_ways_2_mem_port;
  wire                _zz_ways_2_mem_port_1;
  wire       [21:0]   _zz_ways_3_mem_port;
  wire                _zz_ways_3_mem_port_1;
  wire       [3:0]    _zz_status_mem_port;
  wire       [0:0]    _zz_status_loadRead_rsp_0_dirty_1;
  wire       [0:0]    _zz_status_loadRead_rsp_1_dirty;
  wire       [0:0]    _zz_status_loadRead_rsp_2_dirty;
  wire       [0:0]    _zz_status_loadRead_rsp_3_dirty;
  wire       [0:0]    _zz_status_storeRead_rsp_0_dirty_1;
  wire       [0:0]    _zz_status_storeRead_rsp_1_dirty;
  wire       [0:0]    _zz_status_storeRead_rsp_2_dirty;
  wire       [0:0]    _zz_status_storeRead_rsp_3_dirty;
  wire       [1:0]    _zz_wayRandom_valueNext;
  wire       [0:0]    _zz_wayRandom_valueNext_1;
  wire       [2:0]    _zz_plru_ram_port;
  wire       [1:0]    _zz_refill_free_1;
  wire       [1:0]    _zz_refill_free_2;
  reg        [25:0]   _zz_refill_read_cmdAddress;
  reg        [31:0]   _zz_refill_read_rspAddress;
  reg        [1:0]    _zz_refill_read_way;
  wire       [1:0]    _zz_writeback_free_1;
  wire       [1:0]    _zz_writeback_free_2;
  reg        [31:0]   _zz_writeback_read_address;
  reg        [1:0]    _zz_writeback_read_way;
  wire       [2:0]    _zz_writeback_read_wordIndex;
  wire       [0:0]    _zz_writeback_read_wordIndex_1;
  reg        [63:0]   _zz_writeback_read_readedData;
  reg        [31:0]   _zz_writeback_write_bufferRead_payload_address;
  wire       [2:0]    _zz_writeback_write_wordIndex;
  wire       [0:0]    _zz_writeback_write_wordIndex_1;
  reg        [31:0]   _zz_load_pipeline_stages_1_BANKS_MUXES_0;
  wire       [0:0]    _zz_load_pipeline_stages_1_BANKS_MUXES_0_1;
  reg        [31:0]   _zz_load_pipeline_stages_1_BANKS_MUXES_1;
  wire       [0:0]    _zz_load_pipeline_stages_1_BANKS_MUXES_1_1;
  reg        [31:0]   _zz_load_pipeline_stages_1_BANKS_MUXES_2;
  wire       [0:0]    _zz_load_pipeline_stages_1_BANKS_MUXES_2_1;
  reg        [31:0]   _zz_load_pipeline_stages_1_BANKS_MUXES_3;
  wire       [0:0]    _zz_load_pipeline_stages_1_BANKS_MUXES_3_1;
  reg                 _zz__zz_refill_push_payload_victim;
  reg                 _zz_load_ctrl_refillWayNeedWriteback;
  reg        [19:0]   _zz_writeback_push_payload_address;
  reg                 _zz_store_ctrl_replacedWayNeedWriteback;
  reg                 _zz_store_ctrl_replacedWayNeedWriteback_1;
  reg        [19:0]   _zz_writeback_push_payload_address_1;
  reg                 _zz_refill_push_payload_victim_1;
  wire                store_pipeline_stages_0_isThrown;
  wire                store_pipeline_stages_1_isThrown;
  wire                store_pipeline_stages_2_isThrown;
  reg                 store_pipeline_stages_1_FLUSH_FREE;
  reg        [3:0]    store_pipeline_stages_1_CPU_MASK;
  reg        [31:0]   store_pipeline_stages_1_CPU_WORD;
  reg                 store_pipeline_stages_1_IO;
  reg                 store_pipeline_stages_1_FLUSH;
  reg                 store_pipeline_stages_1_PREFETCH;
  reg                 store_pipeline_stages_1_GENERATION;
  reg                 store_pipeline_stages_2_FLUSH_FREE;
  reg        [3:0]    store_pipeline_stages_2_CPU_MASK;
  reg        [31:0]   store_pipeline_stages_2_CPU_WORD;
  reg                 store_pipeline_stages_2_IO;
  wire       [1:0]    store_pipeline_stages_2_REFILL_SLOT;
  wire                store_pipeline_stages_2_REFILL_SLOT_FULL;
  reg                 store_pipeline_stages_2_WAYS_HIT;
  reg                 store_pipeline_stages_2_MISS;
  reg                 store_pipeline_stages_2_REDO;
  reg                 store_pipeline_stages_2_FLUSH;
  wire       [3:0]    store_pipeline_stages_2_WAYS_HAZARD_resulting;
  reg        [3:0]    store_pipeline_stages_2_WAYS_HITS;
  reg                 store_pipeline_stages_2_STATUS_0_dirty;
  reg                 store_pipeline_stages_2_STATUS_1_dirty;
  reg                 store_pipeline_stages_2_STATUS_2_dirty;
  reg                 store_pipeline_stages_2_STATUS_3_dirty;
  reg                 store_pipeline_stages_2_WAYS_TAGS_0_loaded;
  reg        [19:0]   store_pipeline_stages_2_WAYS_TAGS_0_address;
  reg                 store_pipeline_stages_2_WAYS_TAGS_0_fault;
  reg                 store_pipeline_stages_2_WAYS_TAGS_1_loaded;
  reg        [19:0]   store_pipeline_stages_2_WAYS_TAGS_1_address;
  reg                 store_pipeline_stages_2_WAYS_TAGS_1_fault;
  reg                 store_pipeline_stages_2_WAYS_TAGS_2_loaded;
  reg        [19:0]   store_pipeline_stages_2_WAYS_TAGS_2_address;
  reg                 store_pipeline_stages_2_WAYS_TAGS_2_fault;
  reg                 store_pipeline_stages_2_WAYS_TAGS_3_loaded;
  reg        [19:0]   store_pipeline_stages_2_WAYS_TAGS_3_address;
  reg                 store_pipeline_stages_2_WAYS_TAGS_3_fault;
  reg                 store_pipeline_stages_2_PREFETCH;
  reg                 store_pipeline_stages_2_GENERATION;
  wire                store_pipeline_stages_2_GENERATION_OK;
  reg        [0:0]    store_pipeline_stages_2_PLRU_0;
  reg        [1:0]    store_pipeline_stages_2_PLRU_1;
  wire                store_pipeline_stages_2_PROBE;
  reg        [1:0]    store_pipeline_stages_2_REFILL_HITS_EARLY;
  wire       [1:0]    store_pipeline_stages_2_REFILL_HITS;
  reg        [1:0]    store_pipeline_stages_1_REFILL_HITS_EARLY;
  wire                store_pipeline_stages_1_STATUS_overloaded_0_dirty;
  wire                store_pipeline_stages_1_STATUS_overloaded_1_dirty;
  wire                store_pipeline_stages_1_STATUS_overloaded_2_dirty;
  wire                store_pipeline_stages_1_STATUS_overloaded_3_dirty;
  wire                store_pipeline_stages_1_STATUS_0_dirty;
  wire                store_pipeline_stages_1_STATUS_1_dirty;
  wire                store_pipeline_stages_1_STATUS_2_dirty;
  wire                store_pipeline_stages_1_STATUS_3_dirty;
  wire                store_pipeline_stages_1_WAYS_HIT;
  reg        [3:0]    store_pipeline_stages_1_WAYS_HITS;
  wire                store_pipeline_stages_1_WAYS_TAGS_0_loaded;
  wire       [19:0]   store_pipeline_stages_1_WAYS_TAGS_0_address;
  wire                store_pipeline_stages_1_WAYS_TAGS_0_fault;
  wire                store_pipeline_stages_1_WAYS_TAGS_1_loaded;
  wire       [19:0]   store_pipeline_stages_1_WAYS_TAGS_1_address;
  wire                store_pipeline_stages_1_WAYS_TAGS_1_fault;
  wire                store_pipeline_stages_1_WAYS_TAGS_2_loaded;
  wire       [19:0]   store_pipeline_stages_1_WAYS_TAGS_2_address;
  wire                store_pipeline_stages_1_WAYS_TAGS_2_fault;
  wire                store_pipeline_stages_1_WAYS_TAGS_3_loaded;
  wire       [19:0]   store_pipeline_stages_1_WAYS_TAGS_3_address;
  wire                store_pipeline_stages_1_WAYS_TAGS_3_fault;
  wire                store_pipeline_stages_1_ready;
  wire       [0:0]    store_pipeline_stages_1_PLRU_0;
  wire       [1:0]    store_pipeline_stages_1_PLRU_1;
  wire       [3:0]    store_pipeline_stages_0_WAYS_HAZARD;
  wire                store_pipeline_stages_0_GENERATION;
  wire                store_pipeline_stages_0_PREFETCH;
  wire                store_pipeline_stages_0_FLUSH_FREE;
  wire                store_pipeline_stages_0_FLUSH;
  wire                store_pipeline_stages_0_IO;
  wire       [3:0]    store_pipeline_stages_0_CPU_MASK;
  wire       [31:0]   store_pipeline_stages_0_CPU_WORD;
  wire       [31:0]   store_pipeline_stages_0_ADDRESS_POST_TRANSLATION;
  reg        [31:0]   store_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
  reg        [3:0]    store_pipeline_stages_2_WAYS_HAZARD;
  wire       [3:0]    store_pipeline_stages_2_WAYS_HAZARD_overloaded;
  reg        [31:0]   store_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
  reg        [3:0]    store_pipeline_stages_1_WAYS_HAZARD;
  wire       [3:0]    store_pipeline_stages_1_WAYS_HAZARD_overloaded;
  wire                load_pipeline_stages_0_isThrown;
  wire                load_pipeline_stages_1_isThrown;
  wire                load_pipeline_stages_2_isThrown;
  reg                 load_pipeline_stages_1_NEED_UNIQUE;
  wire       [1:0]    load_pipeline_stages_2_REFILL_SLOT;
  wire                load_pipeline_stages_2_REFILL_SLOT_FULL;
  reg                 load_pipeline_stages_2_ABORD;
  wire                load_pipeline_stages_2_FAULT;
  reg                 load_pipeline_stages_2_MISS;
  reg                 load_pipeline_stages_2_LOCKED;
  reg                 load_pipeline_stages_2_REDO;
  reg                 load_pipeline_stages_2_NEED_UNIQUE;
  wire       [3:0]    load_pipeline_stages_2_WAYS_HAZARD_resulting;
  reg        [3:0]    load_pipeline_stages_2_BANK_BUSY_REMAPPED;
  reg                 load_pipeline_stages_2_STATUS_0_dirty;
  reg                 load_pipeline_stages_2_STATUS_1_dirty;
  reg                 load_pipeline_stages_2_STATUS_2_dirty;
  reg                 load_pipeline_stages_2_STATUS_3_dirty;
  reg                 load_pipeline_stages_2_WAYS_TAGS_0_loaded;
  reg        [19:0]   load_pipeline_stages_2_WAYS_TAGS_0_address;
  reg                 load_pipeline_stages_2_WAYS_TAGS_0_fault;
  reg                 load_pipeline_stages_2_WAYS_TAGS_1_loaded;
  reg        [19:0]   load_pipeline_stages_2_WAYS_TAGS_1_address;
  reg                 load_pipeline_stages_2_WAYS_TAGS_1_fault;
  reg                 load_pipeline_stages_2_WAYS_TAGS_2_loaded;
  reg        [19:0]   load_pipeline_stages_2_WAYS_TAGS_2_address;
  reg                 load_pipeline_stages_2_WAYS_TAGS_2_fault;
  reg                 load_pipeline_stages_2_WAYS_TAGS_3_loaded;
  reg        [19:0]   load_pipeline_stages_2_WAYS_TAGS_3_address;
  reg                 load_pipeline_stages_2_WAYS_TAGS_3_fault;
  reg        [0:0]    load_pipeline_stages_2_PLRU_0;
  reg        [1:0]    load_pipeline_stages_2_PLRU_1;
  reg                 load_pipeline_stages_1_UNLOCKED;
  wire                load_pipeline_stages_1_LOCKED;
  reg        [31:0]   load_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
  wire       [1:0]    load_pipeline_stages_2_REFILL_HITS;
  wire                load_pipeline_stages_1_STATUS_overloaded_0_dirty;
  wire                load_pipeline_stages_1_STATUS_overloaded_1_dirty;
  wire                load_pipeline_stages_1_STATUS_overloaded_2_dirty;
  wire                load_pipeline_stages_1_STATUS_overloaded_3_dirty;
  wire                load_pipeline_stages_1_STATUS_0_dirty;
  wire                load_pipeline_stages_1_STATUS_1_dirty;
  wire                load_pipeline_stages_1_STATUS_2_dirty;
  wire                load_pipeline_stages_1_STATUS_3_dirty;
  wire                load_pipeline_stages_2_WAYS_HIT;
  reg        [3:0]    load_pipeline_stages_1_WAYS_HITS;
  wire                load_pipeline_stages_1_WAYS_TAGS_0_loaded;
  wire       [19:0]   load_pipeline_stages_1_WAYS_TAGS_0_address;
  wire                load_pipeline_stages_1_WAYS_TAGS_0_fault;
  wire                load_pipeline_stages_1_WAYS_TAGS_1_loaded;
  wire       [19:0]   load_pipeline_stages_1_WAYS_TAGS_1_address;
  wire                load_pipeline_stages_1_WAYS_TAGS_1_fault;
  wire                load_pipeline_stages_1_WAYS_TAGS_2_loaded;
  wire       [19:0]   load_pipeline_stages_1_WAYS_TAGS_2_address;
  wire                load_pipeline_stages_1_WAYS_TAGS_2_fault;
  wire                load_pipeline_stages_1_WAYS_TAGS_3_loaded;
  wire       [19:0]   load_pipeline_stages_1_WAYS_TAGS_3_address;
  wire                load_pipeline_stages_1_WAYS_TAGS_3_fault;
  wire                load_pipeline_stages_1_ready;
  wire       [0:0]    load_pipeline_stages_1_PLRU_0;
  wire       [1:0]    load_pipeline_stages_1_PLRU_1;
  wire                load_pipeline_stages_1_ABORD;
  wire       [31:0]   load_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
  reg        [31:0]   load_pipeline_stages_2_BANKS_MUXES_0;
  reg        [31:0]   load_pipeline_stages_2_BANKS_MUXES_1;
  reg        [31:0]   load_pipeline_stages_2_BANKS_MUXES_2;
  reg        [31:0]   load_pipeline_stages_2_BANKS_MUXES_3;
  reg        [3:0]    load_pipeline_stages_2_WAYS_HITS;
  wire       [31:0]   load_pipeline_stages_2_CPU_WORD;
  wire       [31:0]   load_pipeline_stages_1_BANKS_MUXES_0;
  wire       [31:0]   load_pipeline_stages_1_BANKS_MUXES_1;
  wire       [31:0]   load_pipeline_stages_1_BANKS_MUXES_2;
  wire       [31:0]   load_pipeline_stages_1_BANKS_MUXES_3;
  reg        [3:0]    load_pipeline_stages_1_BANK_BUSY;
  reg        [3:0]    load_pipeline_stages_1_BANK_BUSY_REMAPPED;
  wire       [63:0]   load_pipeline_stages_1_BANKS_WORDS_0;
  wire       [63:0]   load_pipeline_stages_1_BANKS_WORDS_1;
  wire       [63:0]   load_pipeline_stages_1_BANKS_WORDS_2;
  wire       [63:0]   load_pipeline_stages_1_BANKS_WORDS_3;
  reg        [3:0]    load_pipeline_stages_0_BANK_BUSY_overloaded;
  wire                load_pipeline_stages_0_ready;
  reg        [3:0]    load_pipeline_stages_0_BANK_BUSY;
  wire                load_pipeline_stages_0_NEED_UNIQUE;
  wire                load_pipeline_stages_0_UNLOCKED;
  wire       [3:0]    load_pipeline_stages_0_WAYS_HAZARD;
  wire                load_pipeline_stages_0_REDO_ON_DATA_HAZARD;
  wire       [31:0]   load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION;
  reg        [31:0]   load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION;
  reg        [3:0]    load_pipeline_stages_2_WAYS_HAZARD;
  wire       [3:0]    load_pipeline_stages_2_WAYS_HAZARD_overloaded;
  reg        [31:0]   load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION;
  reg        [3:0]    load_pipeline_stages_1_WAYS_HAZARD;
  wire       [3:0]    load_pipeline_stages_1_WAYS_HAZARD_overloaded;
  reg                 _zz_when_MultiportRam_l328;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 banks_0_write_valid;
  reg        [8:0]    banks_0_write_payload_address;
  reg        [63:0]   banks_0_write_payload_data;
  reg        [7:0]    banks_0_write_payload_mask;
  reg                 banks_0_read_usedByWriteBack;
  reg                 banks_0_read_cmd_valid;
  reg        [8:0]    banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  reg                 banks_1_write_valid;
  reg        [8:0]    banks_1_write_payload_address;
  reg        [63:0]   banks_1_write_payload_data;
  reg        [7:0]    banks_1_write_payload_mask;
  reg                 banks_1_read_usedByWriteBack;
  reg                 banks_1_read_cmd_valid;
  reg        [8:0]    banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  reg                 banks_2_write_valid;
  reg        [8:0]    banks_2_write_payload_address;
  reg        [63:0]   banks_2_write_payload_data;
  reg        [7:0]    banks_2_write_payload_mask;
  reg                 banks_2_read_usedByWriteBack;
  reg                 banks_2_read_cmd_valid;
  reg        [8:0]    banks_2_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   banks_2_read_rsp /* synthesis syn_keep = 1 */ ;
  reg                 banks_3_write_valid;
  reg        [8:0]    banks_3_write_payload_address;
  reg        [63:0]   banks_3_write_payload_data;
  reg        [7:0]    banks_3_write_payload_mask;
  reg                 banks_3_read_usedByWriteBack;
  reg                 banks_3_read_cmd_valid;
  reg        [8:0]    banks_3_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   banks_3_read_rsp /* synthesis syn_keep = 1 */ ;
  reg        [3:0]    waysWrite_mask;
  reg        [5:0]    waysWrite_address;
  reg                 waysWrite_tag_loaded;
  reg        [19:0]   waysWrite_tag_address;
  reg                 waysWrite_tag_fault;
  reg        [3:0]    waysWrite_maskLast;
  reg        [5:0]    waysWrite_addressLast;
  wire                ways_0_loadRead_cmd_valid;
  wire       [5:0]    ways_0_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_0_loadRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   ways_0_loadRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_0_loadRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_ways_0_loadRead_rsp_loaded;
  wire                ways_0_storeRead_cmd_valid;
  wire       [5:0]    ways_0_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_0_storeRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   ways_0_storeRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_0_storeRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_ways_0_storeRead_rsp_loaded;
  wire                ways_1_loadRead_cmd_valid;
  wire       [5:0]    ways_1_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_1_loadRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   ways_1_loadRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_1_loadRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_ways_1_loadRead_rsp_loaded;
  wire                ways_1_storeRead_cmd_valid;
  wire       [5:0]    ways_1_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_1_storeRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   ways_1_storeRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_1_storeRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_ways_1_storeRead_rsp_loaded;
  wire                ways_2_loadRead_cmd_valid;
  wire       [5:0]    ways_2_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_2_loadRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   ways_2_loadRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_2_loadRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_ways_2_loadRead_rsp_loaded;
  wire                ways_2_storeRead_cmd_valid;
  wire       [5:0]    ways_2_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_2_storeRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   ways_2_storeRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_2_storeRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_ways_2_storeRead_rsp_loaded;
  wire                ways_3_loadRead_cmd_valid;
  wire       [5:0]    ways_3_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_3_loadRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   ways_3_loadRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_3_loadRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_ways_3_loadRead_rsp_loaded;
  wire                ways_3_storeRead_cmd_valid;
  wire       [5:0]    ways_3_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                ways_3_storeRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   ways_3_storeRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                ways_3_storeRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_ways_3_storeRead_rsp_loaded;
  reg                 status_write_valid;
  reg        [5:0]    status_write_payload_address;
  reg                 status_write_payload_data_0_dirty;
  reg                 status_write_payload_data_1_dirty;
  reg                 status_write_payload_data_2_dirty;
  reg                 status_write_payload_data_3_dirty;
  wire                status_loadRead_cmd_valid;
  wire       [5:0]    status_loadRead_cmd_payload;
  (* keep , syn_keep *) wire                status_loadRead_rsp_0_dirty /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                status_loadRead_rsp_1_dirty /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                status_loadRead_rsp_2_dirty /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                status_loadRead_rsp_3_dirty /* synthesis syn_keep = 1 */ ;
  wire       [3:0]    _zz_status_loadRead_rsp_0_dirty;
  wire                status_storeRead_cmd_valid;
  wire       [5:0]    status_storeRead_cmd_payload;
  (* keep , syn_keep *) wire                status_storeRead_rsp_0_dirty /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                status_storeRead_rsp_1_dirty /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                status_storeRead_rsp_2_dirty /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                status_storeRead_rsp_3_dirty /* synthesis syn_keep = 1 */ ;
  wire       [3:0]    _zz_status_storeRead_rsp_0_dirty;
  reg                 status_writeLast_valid;
  reg        [5:0]    status_writeLast_payload_address;
  reg                 status_writeLast_payload_data_0_dirty;
  reg                 status_writeLast_payload_data_1_dirty;
  reg                 status_writeLast_payload_data_2_dirty;
  reg                 status_writeLast_payload_data_3_dirty;
  wire                wayRandom_willIncrement;
  wire                wayRandom_willClear;
  reg        [1:0]    wayRandom_valueNext;
  reg        [1:0]    wayRandom_value;
  wire                wayRandom_willOverflowIfInc;
  wire                wayRandom_willOverflow;
  reg                 plru_write_valid;
  reg        [5:0]    plru_write_payload_address;
  reg        [0:0]    plru_write_payload_data_0;
  reg        [1:0]    plru_write_payload_data_1;
  reg                 plru_fromLoad_valid;
  wire       [5:0]    plru_fromLoad_payload_address;
  wire       [0:0]    plru_fromLoad_payload_data_0;
  wire       [1:0]    plru_fromLoad_payload_data_1;
  reg                 plru_fromStore_valid;
  wire       [5:0]    plru_fromStore_payload_address;
  wire       [0:0]    plru_fromStore_payload_data_0;
  wire       [1:0]    plru_fromStore_payload_data_1;
  reg        [6:0]    invalidate_counter;
  wire                invalidate_done;
  wire                invalidate_reservation_win;
  reg                 invalidate_reservation_take;
  wire                when_DataCache_l887;
  reg                 invalidate_firstEver;
  wire                when_DataCache_l896;
  wire       [2:0]    _zz_plru_write_payload_data_0;
  reg                 refill_slots_0_valid;
  reg        [31:0]   refill_slots_0_address;
  reg        [1:0]    refill_slots_0_way;
  reg                 refill_slots_0_cmdSent;
  reg        [0:0]    refill_slots_0_priority;
  reg                 refill_slots_0_loaded;
  reg        [0:0]    refill_slots_0_loadedCounter;
  wire                refill_slots_0_loadedDone;
  wire                when_DataCache_l933;
  wire                refill_slots_0_free;
  reg        [1:0]    refill_slots_0_victim;
  reg        [1:0]    refill_slots_0_writebackHazards;
  reg                 refill_slots_1_valid;
  reg        [31:0]   refill_slots_1_address;
  reg        [1:0]    refill_slots_1_way;
  reg                 refill_slots_1_cmdSent;
  reg        [0:0]    refill_slots_1_priority;
  reg                 refill_slots_1_loaded;
  reg        [0:0]    refill_slots_1_loadedCounter;
  wire                refill_slots_1_loadedDone;
  wire                when_DataCache_l933_1;
  wire                refill_slots_1_free;
  reg        [1:0]    refill_slots_1_victim;
  reg        [1:0]    refill_slots_1_writebackHazards;
  wire       [1:0]    _zz_refill_free;
  wire       [1:0]    refill_free;
  wire                refill_full;
  reg                 refill_push_valid;
  reg        [31:0]   refill_push_payload_address;
  reg        [1:0]    refill_push_payload_way;
  reg        [1:0]    refill_push_payload_victim;
  reg                 refill_push_payload_unique;
  reg                 refill_push_payload_data;
  reg        [31:0]   refill_pushCounter;
  wire                when_DataCache_l960;
  wire                _zz_27;
  wire                _zz_28;
  wire                when_DataCache_l960_1;
  wire                refill_read_arbiter_slotsWithId_0_0;
  wire                refill_read_arbiter_slotsWithId_1_0;
  wire       [1:0]    refill_read_arbiter_hits;
  wire                refill_read_arbiter_hit;
  reg        [1:0]    refill_read_arbiter_oh;
  wire                _zz_refill_read_arbiter_sel;
  wire       [0:0]    refill_read_arbiter_sel;
  reg        [1:0]    refill_read_arbiter_lock;
  wire                when_DataCache_l910;
  reg        [1:0]    refill_read_writebackHazards;
  wire                refill_read_writebackHazard;
  wire                io_mem_read_cmd_fire;
  wire                when_DataCache_l985;
  wire       [31:0]   refill_read_cmdAddress;
  wire                when_DataCache_l997;
  wire                when_DataCache_l997_1;
  wire       [31:0]   refill_read_rspAddress;
  wire       [1:0]    refill_read_way;
  (* keep , syn_keep *) reg        [2:0]    refill_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                refill_read_rspWithData;
  reg        [3:0]    refill_read_bankWriteNotif;
  reg                 refill_read_hadError;
  wire                when_DataCache_l1025;
  reg                 refill_read_fire;
  wire                refill_read_reservation_win;
  reg                 refill_read_reservation_take;
  wire                refill_read_faulty;
  wire                when_DataCache_l1036;
  reg                 writeback_slots_0_fire;
  reg                 writeback_slots_0_valid;
  reg        [31:0]   writeback_slots_0_address;
  reg        [1:0]    writeback_slots_0_way;
  reg        [0:0]    writeback_slots_0_priority;
  reg                 writeback_slots_0_readCmdDone;
  reg                 writeback_slots_0_victimBufferReady;
  reg                 writeback_slots_0_readRspDone;
  reg                 writeback_slots_0_writeCmdDone;
  wire                writeback_slots_0_free;
  reg                 writeback_slots_1_fire;
  reg                 writeback_slots_1_valid;
  reg        [31:0]   writeback_slots_1_address;
  reg        [1:0]    writeback_slots_1_way;
  reg        [0:0]    writeback_slots_1_priority;
  reg                 writeback_slots_1_readCmdDone;
  reg                 writeback_slots_1_victimBufferReady;
  reg                 writeback_slots_1_readRspDone;
  reg                 writeback_slots_1_writeCmdDone;
  wire                writeback_slots_1_free;
  wire       [1:0]    _zz_writeback_free;
  wire       [1:0]    writeback_free;
  wire                writeback_full;
  reg                 writeback_push_valid;
  reg        [31:0]   writeback_push_payload_address;
  reg        [1:0]    writeback_push_payload_way;
  wire                when_DataCache_l1127;
  wire                when_DataCache_l1127_1;
  wire                writeback_read_arbiter_slotsWithId_0_0;
  wire                writeback_read_arbiter_slotsWithId_1_0;
  wire       [1:0]    writeback_read_arbiter_hits;
  wire                writeback_read_arbiter_hit;
  reg        [1:0]    writeback_read_arbiter_oh;
  wire                _zz_writeback_read_arbiter_sel;
  wire       [0:0]    writeback_read_arbiter_sel;
  reg        [1:0]    writeback_read_arbiter_lock;
  wire                when_DataCache_l910_1;
  wire       [31:0]   writeback_read_address;
  wire       [1:0]    writeback_read_way;
  (* keep , syn_keep *) reg        [2:0]    writeback_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                writeback_read_slotRead_valid;
  wire       [0:0]    writeback_read_slotRead_payload_id;
  wire                writeback_read_slotRead_payload_last;
  wire       [2:0]    writeback_read_slotRead_payload_wordIndex;
  wire       [1:0]    writeback_read_slotRead_payload_way;
  wire                when_DataCache_l1174;
  wire                when_DataCache_l1184;
  wire                when_DataCache_l1184_1;
  wire                when_DataCache_l1184_2;
  wire                when_DataCache_l1184_3;
  reg                 writeback_read_slotReadLast_valid;
  reg        [0:0]    writeback_read_slotReadLast_payload_id;
  reg                 writeback_read_slotReadLast_payload_last;
  reg        [2:0]    writeback_read_slotReadLast_payload_wordIndex;
  reg        [1:0]    writeback_read_slotReadLast_payload_way;
  wire       [63:0]   writeback_read_readedData;
  wire       [3:0]    _zz_when_MultiportRam_l328_1;
  wire                writeback_write_arbiter_slotsWithId_0_0;
  wire                writeback_write_arbiter_slotsWithId_1_0;
  wire       [1:0]    writeback_write_arbiter_hits;
  wire                writeback_write_arbiter_hit;
  reg        [1:0]    writeback_write_arbiter_oh;
  wire                _zz_writeback_write_arbiter_sel;
  wire       [0:0]    writeback_write_arbiter_sel;
  reg        [1:0]    writeback_write_arbiter_lock;
  wire                when_DataCache_l910_2;
  (* keep , syn_keep *) reg        [2:0]    writeback_write_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                writeback_write_last;
  wire                writeback_write_bufferRead_valid;
  reg                 writeback_write_bufferRead_ready;
  wire       [0:0]    writeback_write_bufferRead_payload_id;
  wire       [31:0]   writeback_write_bufferRead_payload_address;
  wire                writeback_write_bufferRead_payload_last;
  wire                writeback_write_bufferRead_fire;
  wire                when_DataCache_l1252;
  wire                writeback_write_cmd_valid;
  wire                writeback_write_cmd_ready;
  wire       [0:0]    writeback_write_cmd_payload_id;
  wire       [31:0]   writeback_write_cmd_payload_address;
  wire                writeback_write_cmd_payload_last;
  reg                 writeback_write_bufferRead_rValid;
  reg        [0:0]    writeback_write_bufferRead_rData_id;
  reg        [31:0]   writeback_write_bufferRead_rData_address;
  reg                 writeback_write_bufferRead_rData_last;
  wire                when_Stream_l369;
  wire       [3:0]    _zz_when_MultiportRam_l328_2;
  wire       [63:0]   writeback_write_word;
  wire                load_pipeline_stages_0_valid;
  reg                 _zz_load_pipeline_stages_1_valid;
  reg                 load_pipeline_stages_1_valid;
  reg                 _zz_load_pipeline_stages_2_valid;
  reg                 load_pipeline_stages_2_valid;
  wire                _zz_load_pipeline_stages_0_throwRequest_DataCache_l1301;
  wire                load_pipeline_stages_0_throwRequest_DataCache_l1301;
  wire                _zz_load_pipeline_stages_1_throwRequest_DataCache_l1301;
  wire                load_pipeline_stages_1_throwRequest_DataCache_l1301;
  wire                load_pipeline_stages_2_throwRequest_DataCache_l1301;
  wire                when_DataCache_l1337;
  wire                when_DataCache_l1337_1;
  wire                when_DataCache_l1337_2;
  wire                when_DataCache_l1337_3;
  wire                _zz_load_pipeline_stages_2_CPU_WORD;
  wire                _zz_load_pipeline_stages_2_CPU_WORD_1;
  wire                _zz_load_pipeline_stages_2_CPU_WORD_2;
  wire       [5:0]    _zz_load_pipeline_stages_1_PLRU_0;
  wire       [2:0]    _zz_load_pipeline_stages_1_PLRU_0_1;
  reg                 _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty;
  reg                 _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty;
  reg                 _zz_load_pipeline_stages_1_STATUS_overloaded_2_dirty;
  reg                 _zz_load_pipeline_stages_1_STATUS_overloaded_3_dirty;
  wire                when_DataCache_l859;
  wire                when_DataCache_l862;
  wire       [0:0]    load_ctrl_plruLogic_core_io_context_state_0;
  wire       [1:0]    load_ctrl_plruLogic_core_io_context_state_1;
  wire       [1:0]    load_ctrl_plruLogic_core_io_evict_id;
  reg        [1:0]    load_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    load_ctrl_plruLogic_core_io_update_state_0;
  reg        [1:0]    load_ctrl_plruLogic_core_io_update_state_1;
  wire                load_ctrl_plruLogic_core_evict_sel_0;
  wire                load_ctrl_plruLogic_core_evict_sel_1;
  wire                load_ctrl_plruLogic_core_evict_logic_0_state;
  wire       [0:0]    load_ctrl_plruLogic_core_evict_logic_1_stateSel;
  wire                load_ctrl_plruLogic_core_evict_logic_1_state;
  wire       [0:0]    load_ctrl_plruLogic_core_update_logic_1_sel;
  wire                load_ctrl_reservation_win;
  reg                 load_ctrl_reservation_take;
  wire       [1:0]    load_ctrl_refillWay;
  wire                _zz_refill_push_payload_victim;
  wire                load_ctrl_refillWayNeedWriteback;
  wire                load_ctrl_refillHit;
  wire                load_ctrl_refillLoaded;
  wire                load_ctrl_lineBusy;
  wire                load_ctrl_bankBusy;
  wire                load_ctrl_waysHitHazard;
  wire                load_ctrl_hitUnique;
  wire                load_ctrl_uniqueMiss;
  wire                load_ctrl_canRefill;
  wire                load_ctrl_askRefill;
  reg                 load_ctrl_askUpgrade;
  wire                load_ctrl_startRefill;
  wire                load_ctrl_startUpgrade;
  wire                _zz_load_ctrl_wayId;
  wire                _zz_load_ctrl_wayId_1;
  wire       [1:0]    load_ctrl_wayId;
  wire                when_DataCache_l1471;
  wire       [3:0]    _zz_32;
  wire                when_DataCache_l1512;
  wire                when_Pipeline_l272;
  wire                when_Pipeline_l272_1;
  wire                store_pipeline_stages_0_valid;
  reg                 _zz_store_pipeline_stages_1_valid;
  reg                 store_pipeline_stages_1_valid;
  reg                 _zz_store_pipeline_stages_2_valid;
  reg                 store_pipeline_stages_2_valid;
  wire                store_pipeline_discardAll;
  wire                store_pipeline_stages_0_throwRequest_DataCache_l1551;
  wire                store_pipeline_stages_1_throwRequest_DataCache_l1551;
  wire                store_pipeline_stages_2_throwRequest_DataCache_l1551;
  reg                 store_target;
  wire       [5:0]    _zz_store_pipeline_stages_1_PLRU_0;
  wire       [2:0]    _zz_store_pipeline_stages_1_PLRU_0_1;
  reg                 _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty;
  reg                 _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty;
  reg                 _zz_store_pipeline_stages_1_STATUS_overloaded_2_dirty;
  reg                 _zz_store_pipeline_stages_1_STATUS_overloaded_3_dirty;
  wire                when_DataCache_l859_1;
  wire                when_DataCache_l862_1;
  wire                store_refillCheckEarly_refillPushHit;
  wire       [0:0]    store_ctrl_plruLogic_core_io_context_state_0;
  wire       [1:0]    store_ctrl_plruLogic_core_io_context_state_1;
  wire       [1:0]    store_ctrl_plruLogic_core_io_evict_id;
  reg        [1:0]    store_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    store_ctrl_plruLogic_core_io_update_state_0;
  reg        [1:0]    store_ctrl_plruLogic_core_io_update_state_1;
  wire                store_ctrl_plruLogic_core_evict_sel_0;
  wire                store_ctrl_plruLogic_core_evict_sel_1;
  wire                store_ctrl_plruLogic_core_evict_logic_0_state;
  wire       [0:0]    store_ctrl_plruLogic_core_evict_logic_1_stateSel;
  wire                store_ctrl_plruLogic_core_evict_logic_1_state;
  wire       [0:0]    store_ctrl_plruLogic_core_update_logic_1_sel;
  wire                store_ctrl_reservation_win;
  reg                 store_ctrl_reservation_take;
  wire       [1:0]    store_ctrl_replacedWay;
  wire                store_ctrl_replacedWayNeedWriteback;
  wire                store_ctrl_refillHit;
  wire                store_ctrl_lineBusy;
  wire                store_ctrl_waysHitHazard;
  wire                store_ctrl_wasClean;
  wire                store_ctrl_bankBusy;
  wire                store_ctrl_hitUnique;
  wire                store_ctrl_hitFault;
  reg        [1:0]    store_ctrl_refillWay;
  wire                store_ctrl_canRefill;
  wire                store_ctrl_askRefill;
  wire                store_ctrl_askUpgrade;
  reg                 store_ctrl_startRefill;
  reg                 store_ctrl_startUpgrade;
  reg                 store_ctrl_writeCache;
  reg                 store_ctrl_setDirty;
  wire                _zz_store_ctrl_wayId;
  wire                _zz_store_ctrl_wayId_1;
  wire                _zz_store_ctrl_wayId_2;
  wire                _zz_store_ctrl_wayId_3;
  wire                _zz_store_ctrl_wayId_4;
  wire       [1:0]    store_ctrl_wayId;
  wire       [3:0]    store_ctrl_needFlushs;
  wire       [3:0]    _zz_store_ctrl_needFlushs_bools_0;
  wire                store_ctrl_needFlushs_bools_0;
  wire                store_ctrl_needFlushs_bools_1;
  wire                store_ctrl_needFlushs_bools_2;
  wire                store_ctrl_needFlushs_bools_3;
  reg        [3:0]    _zz_store_ctrl_needFlushOh;
  wire                store_ctrl_needFlushs_range_0_to_1;
  wire                store_ctrl_needFlushs_range_0_to_2;
  wire       [3:0]    store_ctrl_needFlushOh;
  wire                _zz_34;
  wire                _zz_store_ctrl_needFlushSel;
  wire                _zz_store_ctrl_needFlushSel_1;
  wire                _zz_store_ctrl_needFlushSel_2;
  wire                _zz_store_ctrl_needFlushSel_3;
  wire                _zz_store_ctrl_needFlushSel_4;
  wire       [1:0]    store_ctrl_needFlushSel;
  wire                store_ctrl_needFlush;
  wire                store_ctrl_canFlush;
  wire                store_ctrl_startFlush;
  wire                when_DataCache_l1705;
  wire                when_DataCache_l1725;
  wire                when_DataCache_l1732;
  wire                when_DataCache_l1750;
  wire                when_DataCache_l1774;
  wire       [1:0]    _zz_35;
  wire                when_DataCache_l1774_1;
  wire       [1:0]    _zz_36;
  wire                when_DataCache_l1774_2;
  wire       [1:0]    _zz_37;
  wire                when_DataCache_l1774_3;
  wire       [1:0]    _zz_38;
  wire                when_DataCache_l1804;
  wire                when_Pipeline_l272_2;
  wire                when_Pipeline_l272_3;
  reg        [63:0]   _zz_banks_0_read_rsp;
  reg                 when_MultiportRam_l328;
  reg        [7:0]    _zz_39;
  reg        [63:0]   _zz_banks_1_read_rsp;
  reg                 when_MultiportRam_l328_1;
  reg        [7:0]    _zz_40;
  reg        [63:0]   _zz_banks_2_read_rsp;
  reg                 when_MultiportRam_l328_2;
  reg        [7:0]    _zz_41;
  reg        [63:0]   _zz_banks_3_read_rsp;
  reg                 when_MultiportRam_l328_3;
  reg        [7:0]    _zz_42;
  reg        [63:0]   _zz_writeback_write_word;
  reg                 when_MultiportRam_l328_4;
  reg [7:0] banks_0_mem_symbol0 [0:511];
  reg [7:0] banks_0_mem_symbol1 [0:511];
  reg [7:0] banks_0_mem_symbol2 [0:511];
  reg [7:0] banks_0_mem_symbol3 [0:511];
  reg [7:0] banks_0_mem_symbol4 [0:511];
  reg [7:0] banks_0_mem_symbol5 [0:511];
  reg [7:0] banks_0_mem_symbol6 [0:511];
  reg [7:0] banks_0_mem_symbol7 [0:511];
  reg [7:0] _zz_banks_0_memsymbol_read;
  reg [7:0] _zz_banks_0_memsymbol_read_1;
  reg [7:0] _zz_banks_0_memsymbol_read_2;
  reg [7:0] _zz_banks_0_memsymbol_read_3;
  reg [7:0] _zz_banks_0_memsymbol_read_4;
  reg [7:0] _zz_banks_0_memsymbol_read_5;
  reg [7:0] _zz_banks_0_memsymbol_read_6;
  reg [7:0] _zz_banks_0_memsymbol_read_7;
  reg [7:0] banks_1_mem_symbol0 [0:511];
  reg [7:0] banks_1_mem_symbol1 [0:511];
  reg [7:0] banks_1_mem_symbol2 [0:511];
  reg [7:0] banks_1_mem_symbol3 [0:511];
  reg [7:0] banks_1_mem_symbol4 [0:511];
  reg [7:0] banks_1_mem_symbol5 [0:511];
  reg [7:0] banks_1_mem_symbol6 [0:511];
  reg [7:0] banks_1_mem_symbol7 [0:511];
  reg [7:0] _zz_banks_1_memsymbol_read;
  reg [7:0] _zz_banks_1_memsymbol_read_1;
  reg [7:0] _zz_banks_1_memsymbol_read_2;
  reg [7:0] _zz_banks_1_memsymbol_read_3;
  reg [7:0] _zz_banks_1_memsymbol_read_4;
  reg [7:0] _zz_banks_1_memsymbol_read_5;
  reg [7:0] _zz_banks_1_memsymbol_read_6;
  reg [7:0] _zz_banks_1_memsymbol_read_7;
  reg [7:0] banks_2_mem_symbol0 [0:511];
  reg [7:0] banks_2_mem_symbol1 [0:511];
  reg [7:0] banks_2_mem_symbol2 [0:511];
  reg [7:0] banks_2_mem_symbol3 [0:511];
  reg [7:0] banks_2_mem_symbol4 [0:511];
  reg [7:0] banks_2_mem_symbol5 [0:511];
  reg [7:0] banks_2_mem_symbol6 [0:511];
  reg [7:0] banks_2_mem_symbol7 [0:511];
  reg [7:0] _zz_banks_2_memsymbol_read;
  reg [7:0] _zz_banks_2_memsymbol_read_1;
  reg [7:0] _zz_banks_2_memsymbol_read_2;
  reg [7:0] _zz_banks_2_memsymbol_read_3;
  reg [7:0] _zz_banks_2_memsymbol_read_4;
  reg [7:0] _zz_banks_2_memsymbol_read_5;
  reg [7:0] _zz_banks_2_memsymbol_read_6;
  reg [7:0] _zz_banks_2_memsymbol_read_7;
  reg [7:0] banks_3_mem_symbol0 [0:511];
  reg [7:0] banks_3_mem_symbol1 [0:511];
  reg [7:0] banks_3_mem_symbol2 [0:511];
  reg [7:0] banks_3_mem_symbol3 [0:511];
  reg [7:0] banks_3_mem_symbol4 [0:511];
  reg [7:0] banks_3_mem_symbol5 [0:511];
  reg [7:0] banks_3_mem_symbol6 [0:511];
  reg [7:0] banks_3_mem_symbol7 [0:511];
  reg [7:0] _zz_banks_3_memsymbol_read;
  reg [7:0] _zz_banks_3_memsymbol_read_1;
  reg [7:0] _zz_banks_3_memsymbol_read_2;
  reg [7:0] _zz_banks_3_memsymbol_read_3;
  reg [7:0] _zz_banks_3_memsymbol_read_4;
  reg [7:0] _zz_banks_3_memsymbol_read_5;
  reg [7:0] _zz_banks_3_memsymbol_read_6;
  reg [7:0] _zz_banks_3_memsymbol_read_7;
  (* ram_style = "distributed" *) reg [21:0] ways_0_mem [0:63];
  (* ram_style = "distributed" *) reg [21:0] ways_1_mem [0:63];
  (* ram_style = "distributed" *) reg [21:0] ways_2_mem [0:63];
  (* ram_style = "distributed" *) reg [21:0] ways_3_mem [0:63];
  (* ram_style = "distributed" *) reg [3:0] status_mem [0:63];
  (* ram_style = "distributed" *) reg [2:0] plru_ram [0:63];
  reg [63:0] writeback_victimBuffer [0:15];

  assign _zz_status_loadRead_rsp_0_dirty_1 = _zz_status_loadRead_rsp_0_dirty[0 : 0];
  assign _zz_status_loadRead_rsp_1_dirty = _zz_status_loadRead_rsp_0_dirty[1 : 1];
  assign _zz_status_loadRead_rsp_2_dirty = _zz_status_loadRead_rsp_0_dirty[2 : 2];
  assign _zz_status_loadRead_rsp_3_dirty = _zz_status_loadRead_rsp_0_dirty[3 : 3];
  assign _zz_status_storeRead_rsp_0_dirty_1 = _zz_status_storeRead_rsp_0_dirty[0 : 0];
  assign _zz_status_storeRead_rsp_1_dirty = _zz_status_storeRead_rsp_0_dirty[1 : 1];
  assign _zz_status_storeRead_rsp_2_dirty = _zz_status_storeRead_rsp_0_dirty[2 : 2];
  assign _zz_status_storeRead_rsp_3_dirty = _zz_status_storeRead_rsp_0_dirty[3 : 3];
  assign _zz_wayRandom_valueNext_1 = wayRandom_willIncrement;
  assign _zz_wayRandom_valueNext = {1'd0, _zz_wayRandom_valueNext_1};
  assign _zz_refill_free_1 = (_zz_refill_free & (~ _zz_refill_free_2));
  assign _zz_refill_free_2 = (_zz_refill_free - 2'b01);
  assign _zz_writeback_free_1 = (_zz_writeback_free & (~ _zz_writeback_free_2));
  assign _zz_writeback_free_2 = (_zz_writeback_free - 2'b01);
  assign _zz_writeback_read_wordIndex_1 = writeback_read_slotRead_valid;
  assign _zz_writeback_read_wordIndex = {2'd0, _zz_writeback_read_wordIndex_1};
  assign _zz_writeback_write_wordIndex_1 = (writeback_write_bufferRead_fire && 1'b1);
  assign _zz_writeback_write_wordIndex = {2'd0, _zz_writeback_write_wordIndex_1};
  assign _zz_ways_0_mem_port = {waysWrite_tag_fault,{waysWrite_tag_address,waysWrite_tag_loaded}};
  assign _zz_ways_0_mem_port_1 = waysWrite_mask[0];
  assign _zz_ways_1_mem_port = {waysWrite_tag_fault,{waysWrite_tag_address,waysWrite_tag_loaded}};
  assign _zz_ways_1_mem_port_1 = waysWrite_mask[1];
  assign _zz_ways_2_mem_port = {waysWrite_tag_fault,{waysWrite_tag_address,waysWrite_tag_loaded}};
  assign _zz_ways_2_mem_port_1 = waysWrite_mask[2];
  assign _zz_ways_3_mem_port = {waysWrite_tag_fault,{waysWrite_tag_address,waysWrite_tag_loaded}};
  assign _zz_ways_3_mem_port_1 = waysWrite_mask[3];
  assign _zz_status_mem_port = {status_write_payload_data_3_dirty,{status_write_payload_data_2_dirty,{status_write_payload_data_1_dirty,status_write_payload_data_0_dirty}}};
  assign _zz_plru_ram_port = {plru_write_payload_data_1,plru_write_payload_data_0};
  assign _zz_load_pipeline_stages_1_BANKS_MUXES_0_1 = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[2 : 2];
  assign _zz_load_pipeline_stages_1_BANKS_MUXES_1_1 = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[2 : 2];
  assign _zz_load_pipeline_stages_1_BANKS_MUXES_2_1 = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[2 : 2];
  assign _zz_load_pipeline_stages_1_BANKS_MUXES_3_1 = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[2 : 2];
  always @(*) begin
    _zz_banks_0_mem_port1 = {_zz_banks_0_memsymbol_read_7, _zz_banks_0_memsymbol_read_6, _zz_banks_0_memsymbol_read_5, _zz_banks_0_memsymbol_read_4, _zz_banks_0_memsymbol_read_3, _zz_banks_0_memsymbol_read_2, _zz_banks_0_memsymbol_read_1, _zz_banks_0_memsymbol_read};
  end
  always @(posedge clk) begin
    if(banks_0_write_payload_mask[0] && banks_0_write_valid) begin
      banks_0_mem_symbol0[banks_0_write_payload_address] <= banks_0_write_payload_data[7 : 0];
    end
    if(banks_0_write_payload_mask[1] && banks_0_write_valid) begin
      banks_0_mem_symbol1[banks_0_write_payload_address] <= banks_0_write_payload_data[15 : 8];
    end
    if(banks_0_write_payload_mask[2] && banks_0_write_valid) begin
      banks_0_mem_symbol2[banks_0_write_payload_address] <= banks_0_write_payload_data[23 : 16];
    end
    if(banks_0_write_payload_mask[3] && banks_0_write_valid) begin
      banks_0_mem_symbol3[banks_0_write_payload_address] <= banks_0_write_payload_data[31 : 24];
    end
    if(banks_0_write_payload_mask[4] && banks_0_write_valid) begin
      banks_0_mem_symbol4[banks_0_write_payload_address] <= banks_0_write_payload_data[39 : 32];
    end
    if(banks_0_write_payload_mask[5] && banks_0_write_valid) begin
      banks_0_mem_symbol5[banks_0_write_payload_address] <= banks_0_write_payload_data[47 : 40];
    end
    if(banks_0_write_payload_mask[6] && banks_0_write_valid) begin
      banks_0_mem_symbol6[banks_0_write_payload_address] <= banks_0_write_payload_data[55 : 48];
    end
    if(banks_0_write_payload_mask[7] && banks_0_write_valid) begin
      banks_0_mem_symbol7[banks_0_write_payload_address] <= banks_0_write_payload_data[63 : 56];
    end
  end

  always @(posedge clk) begin
    if(banks_0_read_cmd_valid) begin
      _zz_banks_0_memsymbol_read <= banks_0_mem_symbol0[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_1 <= banks_0_mem_symbol1[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_2 <= banks_0_mem_symbol2[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_3 <= banks_0_mem_symbol3[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_4 <= banks_0_mem_symbol4[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_5 <= banks_0_mem_symbol5[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_6 <= banks_0_mem_symbol6[banks_0_read_cmd_payload];
      _zz_banks_0_memsymbol_read_7 <= banks_0_mem_symbol7[banks_0_read_cmd_payload];
    end
  end

  always @(*) begin
    _zz_banks_1_mem_port1 = {_zz_banks_1_memsymbol_read_7, _zz_banks_1_memsymbol_read_6, _zz_banks_1_memsymbol_read_5, _zz_banks_1_memsymbol_read_4, _zz_banks_1_memsymbol_read_3, _zz_banks_1_memsymbol_read_2, _zz_banks_1_memsymbol_read_1, _zz_banks_1_memsymbol_read};
  end
  always @(posedge clk) begin
    if(banks_1_write_payload_mask[0] && banks_1_write_valid) begin
      banks_1_mem_symbol0[banks_1_write_payload_address] <= banks_1_write_payload_data[7 : 0];
    end
    if(banks_1_write_payload_mask[1] && banks_1_write_valid) begin
      banks_1_mem_symbol1[banks_1_write_payload_address] <= banks_1_write_payload_data[15 : 8];
    end
    if(banks_1_write_payload_mask[2] && banks_1_write_valid) begin
      banks_1_mem_symbol2[banks_1_write_payload_address] <= banks_1_write_payload_data[23 : 16];
    end
    if(banks_1_write_payload_mask[3] && banks_1_write_valid) begin
      banks_1_mem_symbol3[banks_1_write_payload_address] <= banks_1_write_payload_data[31 : 24];
    end
    if(banks_1_write_payload_mask[4] && banks_1_write_valid) begin
      banks_1_mem_symbol4[banks_1_write_payload_address] <= banks_1_write_payload_data[39 : 32];
    end
    if(banks_1_write_payload_mask[5] && banks_1_write_valid) begin
      banks_1_mem_symbol5[banks_1_write_payload_address] <= banks_1_write_payload_data[47 : 40];
    end
    if(banks_1_write_payload_mask[6] && banks_1_write_valid) begin
      banks_1_mem_symbol6[banks_1_write_payload_address] <= banks_1_write_payload_data[55 : 48];
    end
    if(banks_1_write_payload_mask[7] && banks_1_write_valid) begin
      banks_1_mem_symbol7[banks_1_write_payload_address] <= banks_1_write_payload_data[63 : 56];
    end
  end

  always @(posedge clk) begin
    if(banks_1_read_cmd_valid) begin
      _zz_banks_1_memsymbol_read <= banks_1_mem_symbol0[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_1 <= banks_1_mem_symbol1[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_2 <= banks_1_mem_symbol2[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_3 <= banks_1_mem_symbol3[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_4 <= banks_1_mem_symbol4[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_5 <= banks_1_mem_symbol5[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_6 <= banks_1_mem_symbol6[banks_1_read_cmd_payload];
      _zz_banks_1_memsymbol_read_7 <= banks_1_mem_symbol7[banks_1_read_cmd_payload];
    end
  end

  always @(*) begin
    _zz_banks_2_mem_port1 = {_zz_banks_2_memsymbol_read_7, _zz_banks_2_memsymbol_read_6, _zz_banks_2_memsymbol_read_5, _zz_banks_2_memsymbol_read_4, _zz_banks_2_memsymbol_read_3, _zz_banks_2_memsymbol_read_2, _zz_banks_2_memsymbol_read_1, _zz_banks_2_memsymbol_read};
  end
  always @(posedge clk) begin
    if(banks_2_write_payload_mask[0] && banks_2_write_valid) begin
      banks_2_mem_symbol0[banks_2_write_payload_address] <= banks_2_write_payload_data[7 : 0];
    end
    if(banks_2_write_payload_mask[1] && banks_2_write_valid) begin
      banks_2_mem_symbol1[banks_2_write_payload_address] <= banks_2_write_payload_data[15 : 8];
    end
    if(banks_2_write_payload_mask[2] && banks_2_write_valid) begin
      banks_2_mem_symbol2[banks_2_write_payload_address] <= banks_2_write_payload_data[23 : 16];
    end
    if(banks_2_write_payload_mask[3] && banks_2_write_valid) begin
      banks_2_mem_symbol3[banks_2_write_payload_address] <= banks_2_write_payload_data[31 : 24];
    end
    if(banks_2_write_payload_mask[4] && banks_2_write_valid) begin
      banks_2_mem_symbol4[banks_2_write_payload_address] <= banks_2_write_payload_data[39 : 32];
    end
    if(banks_2_write_payload_mask[5] && banks_2_write_valid) begin
      banks_2_mem_symbol5[banks_2_write_payload_address] <= banks_2_write_payload_data[47 : 40];
    end
    if(banks_2_write_payload_mask[6] && banks_2_write_valid) begin
      banks_2_mem_symbol6[banks_2_write_payload_address] <= banks_2_write_payload_data[55 : 48];
    end
    if(banks_2_write_payload_mask[7] && banks_2_write_valid) begin
      banks_2_mem_symbol7[banks_2_write_payload_address] <= banks_2_write_payload_data[63 : 56];
    end
  end

  always @(posedge clk) begin
    if(banks_2_read_cmd_valid) begin
      _zz_banks_2_memsymbol_read <= banks_2_mem_symbol0[banks_2_read_cmd_payload];
      _zz_banks_2_memsymbol_read_1 <= banks_2_mem_symbol1[banks_2_read_cmd_payload];
      _zz_banks_2_memsymbol_read_2 <= banks_2_mem_symbol2[banks_2_read_cmd_payload];
      _zz_banks_2_memsymbol_read_3 <= banks_2_mem_symbol3[banks_2_read_cmd_payload];
      _zz_banks_2_memsymbol_read_4 <= banks_2_mem_symbol4[banks_2_read_cmd_payload];
      _zz_banks_2_memsymbol_read_5 <= banks_2_mem_symbol5[banks_2_read_cmd_payload];
      _zz_banks_2_memsymbol_read_6 <= banks_2_mem_symbol6[banks_2_read_cmd_payload];
      _zz_banks_2_memsymbol_read_7 <= banks_2_mem_symbol7[banks_2_read_cmd_payload];
    end
  end

  always @(*) begin
    _zz_banks_3_mem_port1 = {_zz_banks_3_memsymbol_read_7, _zz_banks_3_memsymbol_read_6, _zz_banks_3_memsymbol_read_5, _zz_banks_3_memsymbol_read_4, _zz_banks_3_memsymbol_read_3, _zz_banks_3_memsymbol_read_2, _zz_banks_3_memsymbol_read_1, _zz_banks_3_memsymbol_read};
  end
  always @(posedge clk) begin
    if(banks_3_write_payload_mask[0] && banks_3_write_valid) begin
      banks_3_mem_symbol0[banks_3_write_payload_address] <= banks_3_write_payload_data[7 : 0];
    end
    if(banks_3_write_payload_mask[1] && banks_3_write_valid) begin
      banks_3_mem_symbol1[banks_3_write_payload_address] <= banks_3_write_payload_data[15 : 8];
    end
    if(banks_3_write_payload_mask[2] && banks_3_write_valid) begin
      banks_3_mem_symbol2[banks_3_write_payload_address] <= banks_3_write_payload_data[23 : 16];
    end
    if(banks_3_write_payload_mask[3] && banks_3_write_valid) begin
      banks_3_mem_symbol3[banks_3_write_payload_address] <= banks_3_write_payload_data[31 : 24];
    end
    if(banks_3_write_payload_mask[4] && banks_3_write_valid) begin
      banks_3_mem_symbol4[banks_3_write_payload_address] <= banks_3_write_payload_data[39 : 32];
    end
    if(banks_3_write_payload_mask[5] && banks_3_write_valid) begin
      banks_3_mem_symbol5[banks_3_write_payload_address] <= banks_3_write_payload_data[47 : 40];
    end
    if(banks_3_write_payload_mask[6] && banks_3_write_valid) begin
      banks_3_mem_symbol6[banks_3_write_payload_address] <= banks_3_write_payload_data[55 : 48];
    end
    if(banks_3_write_payload_mask[7] && banks_3_write_valid) begin
      banks_3_mem_symbol7[banks_3_write_payload_address] <= banks_3_write_payload_data[63 : 56];
    end
  end

  always @(posedge clk) begin
    if(banks_3_read_cmd_valid) begin
      _zz_banks_3_memsymbol_read <= banks_3_mem_symbol0[banks_3_read_cmd_payload];
      _zz_banks_3_memsymbol_read_1 <= banks_3_mem_symbol1[banks_3_read_cmd_payload];
      _zz_banks_3_memsymbol_read_2 <= banks_3_mem_symbol2[banks_3_read_cmd_payload];
      _zz_banks_3_memsymbol_read_3 <= banks_3_mem_symbol3[banks_3_read_cmd_payload];
      _zz_banks_3_memsymbol_read_4 <= banks_3_mem_symbol4[banks_3_read_cmd_payload];
      _zz_banks_3_memsymbol_read_5 <= banks_3_mem_symbol5[banks_3_read_cmd_payload];
      _zz_banks_3_memsymbol_read_6 <= banks_3_mem_symbol6[banks_3_read_cmd_payload];
      _zz_banks_3_memsymbol_read_7 <= banks_3_mem_symbol7[banks_3_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_ways_0_mem_port_1) begin
      ways_0_mem[waysWrite_address] <= _zz_ways_0_mem_port;
    end
  end

  assign _zz_ways_0_mem_port1 = ways_0_mem[ways_0_loadRead_cmd_payload];
  assign _zz_ways_0_mem_port2 = ways_0_mem[ways_0_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_ways_1_mem_port_1) begin
      ways_1_mem[waysWrite_address] <= _zz_ways_1_mem_port;
    end
  end

  assign _zz_ways_1_mem_port1 = ways_1_mem[ways_1_loadRead_cmd_payload];
  assign _zz_ways_1_mem_port2 = ways_1_mem[ways_1_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_ways_2_mem_port_1) begin
      ways_2_mem[waysWrite_address] <= _zz_ways_2_mem_port;
    end
  end

  assign _zz_ways_2_mem_port1 = ways_2_mem[ways_2_loadRead_cmd_payload];
  assign _zz_ways_2_mem_port2 = ways_2_mem[ways_2_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_ways_3_mem_port_1) begin
      ways_3_mem[waysWrite_address] <= _zz_ways_3_mem_port;
    end
  end

  assign _zz_ways_3_mem_port1 = ways_3_mem[ways_3_loadRead_cmd_payload];
  assign _zz_ways_3_mem_port2 = ways_3_mem[ways_3_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_2) begin
      status_mem[status_write_payload_address] <= _zz_status_mem_port;
    end
  end

  assign _zz_status_mem_port1 = status_mem[status_loadRead_cmd_payload];
  assign _zz_status_mem_port2 = status_mem[status_storeRead_cmd_payload];
  always @(posedge clk) begin
    if(_zz_1) begin
      plru_ram[plru_write_payload_address] <= _zz_plru_ram_port;
    end
  end

  assign _zz_plru_ram_port1 = plru_ram[_zz_load_pipeline_stages_1_PLRU_0];
  assign _zz_plru_ram_port2 = plru_ram[_zz_store_pipeline_stages_1_PLRU_0];
  always @(posedge clk) begin
    if(_zz_when_MultiportRam_l328) begin
      writeback_victimBuffer[_zz_when_MultiportRam_l328_1] <= writeback_read_readedData;
    end
  end

  always @(posedge clk) begin
    if(writeback_write_bufferRead_ready) begin
      _zz_writeback_victimBuffer_port1 <= writeback_victimBuffer[_zz_when_MultiportRam_l328_2];
    end
  end

  always @(*) begin
    case(refill_read_arbiter_sel)
      1'b0 : _zz_refill_read_cmdAddress = refill_slots_0_address[31 : 6];
      default : _zz_refill_read_cmdAddress = refill_slots_1_address[31 : 6];
    endcase
  end

  always @(*) begin
    case(io_mem_read_rsp_payload_id)
      1'b0 : begin
        _zz_refill_read_rspAddress = refill_slots_0_address;
        _zz_refill_read_way = refill_slots_0_way;
      end
      default : begin
        _zz_refill_read_rspAddress = refill_slots_1_address;
        _zz_refill_read_way = refill_slots_1_way;
      end
    endcase
  end

  always @(*) begin
    case(writeback_read_arbiter_sel)
      1'b0 : begin
        _zz_writeback_read_address = writeback_slots_0_address;
        _zz_writeback_read_way = writeback_slots_0_way;
      end
      default : begin
        _zz_writeback_read_address = writeback_slots_1_address;
        _zz_writeback_read_way = writeback_slots_1_way;
      end
    endcase
  end

  always @(*) begin
    case(writeback_read_slotReadLast_payload_way)
      2'b00 : _zz_writeback_read_readedData = banks_0_read_rsp;
      2'b01 : _zz_writeback_read_readedData = banks_1_read_rsp;
      2'b10 : _zz_writeback_read_readedData = banks_2_read_rsp;
      default : _zz_writeback_read_readedData = banks_3_read_rsp;
    endcase
  end

  always @(*) begin
    case(writeback_write_arbiter_sel)
      1'b0 : _zz_writeback_write_bufferRead_payload_address = writeback_slots_0_address;
      default : _zz_writeback_write_bufferRead_payload_address = writeback_slots_1_address;
    endcase
  end

  always @(*) begin
    case(_zz_load_pipeline_stages_1_BANKS_MUXES_0_1)
      1'b0 : _zz_load_pipeline_stages_1_BANKS_MUXES_0 = load_pipeline_stages_1_BANKS_WORDS_0[31 : 0];
      default : _zz_load_pipeline_stages_1_BANKS_MUXES_0 = load_pipeline_stages_1_BANKS_WORDS_0[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_load_pipeline_stages_1_BANKS_MUXES_1_1)
      1'b0 : _zz_load_pipeline_stages_1_BANKS_MUXES_1 = load_pipeline_stages_1_BANKS_WORDS_1[31 : 0];
      default : _zz_load_pipeline_stages_1_BANKS_MUXES_1 = load_pipeline_stages_1_BANKS_WORDS_1[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_load_pipeline_stages_1_BANKS_MUXES_2_1)
      1'b0 : _zz_load_pipeline_stages_1_BANKS_MUXES_2 = load_pipeline_stages_1_BANKS_WORDS_2[31 : 0];
      default : _zz_load_pipeline_stages_1_BANKS_MUXES_2 = load_pipeline_stages_1_BANKS_WORDS_2[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_load_pipeline_stages_1_BANKS_MUXES_3_1)
      1'b0 : _zz_load_pipeline_stages_1_BANKS_MUXES_3 = load_pipeline_stages_1_BANKS_WORDS_3[31 : 0];
      default : _zz_load_pipeline_stages_1_BANKS_MUXES_3 = load_pipeline_stages_1_BANKS_WORDS_3[63 : 32];
    endcase
  end

  always @(*) begin
    case(load_ctrl_refillWay)
      2'b00 : begin
        _zz__zz_refill_push_payload_victim = load_pipeline_stages_2_STATUS_0_dirty;
        _zz_load_ctrl_refillWayNeedWriteback = load_pipeline_stages_2_WAYS_TAGS_0_loaded;
        _zz_writeback_push_payload_address = load_pipeline_stages_2_WAYS_TAGS_0_address;
      end
      2'b01 : begin
        _zz__zz_refill_push_payload_victim = load_pipeline_stages_2_STATUS_1_dirty;
        _zz_load_ctrl_refillWayNeedWriteback = load_pipeline_stages_2_WAYS_TAGS_1_loaded;
        _zz_writeback_push_payload_address = load_pipeline_stages_2_WAYS_TAGS_1_address;
      end
      2'b10 : begin
        _zz__zz_refill_push_payload_victim = load_pipeline_stages_2_STATUS_2_dirty;
        _zz_load_ctrl_refillWayNeedWriteback = load_pipeline_stages_2_WAYS_TAGS_2_loaded;
        _zz_writeback_push_payload_address = load_pipeline_stages_2_WAYS_TAGS_2_address;
      end
      default : begin
        _zz__zz_refill_push_payload_victim = load_pipeline_stages_2_STATUS_3_dirty;
        _zz_load_ctrl_refillWayNeedWriteback = load_pipeline_stages_2_WAYS_TAGS_3_loaded;
        _zz_writeback_push_payload_address = load_pipeline_stages_2_WAYS_TAGS_3_address;
      end
    endcase
  end

  always @(*) begin
    case(store_ctrl_replacedWay)
      2'b00 : begin
        _zz_store_ctrl_replacedWayNeedWriteback = store_pipeline_stages_2_WAYS_TAGS_0_loaded;
        _zz_store_ctrl_replacedWayNeedWriteback_1 = store_pipeline_stages_2_STATUS_0_dirty;
      end
      2'b01 : begin
        _zz_store_ctrl_replacedWayNeedWriteback = store_pipeline_stages_2_WAYS_TAGS_1_loaded;
        _zz_store_ctrl_replacedWayNeedWriteback_1 = store_pipeline_stages_2_STATUS_1_dirty;
      end
      2'b10 : begin
        _zz_store_ctrl_replacedWayNeedWriteback = store_pipeline_stages_2_WAYS_TAGS_2_loaded;
        _zz_store_ctrl_replacedWayNeedWriteback_1 = store_pipeline_stages_2_STATUS_2_dirty;
      end
      default : begin
        _zz_store_ctrl_replacedWayNeedWriteback = store_pipeline_stages_2_WAYS_TAGS_3_loaded;
        _zz_store_ctrl_replacedWayNeedWriteback_1 = store_pipeline_stages_2_STATUS_3_dirty;
      end
    endcase
  end

  always @(*) begin
    case(writeback_push_payload_way)
      2'b00 : _zz_writeback_push_payload_address_1 = store_pipeline_stages_2_WAYS_TAGS_0_address;
      2'b01 : _zz_writeback_push_payload_address_1 = store_pipeline_stages_2_WAYS_TAGS_1_address;
      2'b10 : _zz_writeback_push_payload_address_1 = store_pipeline_stages_2_WAYS_TAGS_2_address;
      default : _zz_writeback_push_payload_address_1 = store_pipeline_stages_2_WAYS_TAGS_3_address;
    endcase
  end

  always @(*) begin
    case(store_ctrl_refillWay)
      2'b00 : _zz_refill_push_payload_victim_1 = store_pipeline_stages_2_STATUS_0_dirty;
      2'b01 : _zz_refill_push_payload_victim_1 = store_pipeline_stages_2_STATUS_1_dirty;
      2'b10 : _zz_refill_push_payload_victim_1 = store_pipeline_stages_2_STATUS_2_dirty;
      default : _zz_refill_push_payload_victim_1 = store_pipeline_stages_2_STATUS_3_dirty;
    endcase
  end

  always @(*) begin
    _zz_when_MultiportRam_l328 = 1'b0;
    if(writeback_read_slotReadLast_valid) begin
      _zz_when_MultiportRam_l328 = 1'b1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(plru_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(status_write_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    banks_0_read_usedByWriteBack = 1'b0;
    if(when_DataCache_l1184) begin
      banks_0_read_usedByWriteBack = 1'b1;
    end
  end

  assign banks_0_read_rsp = _zz_banks_0_read_rsp;
  always @(*) begin
    banks_0_read_cmd_valid = 1'b0;
    if(when_DataCache_l1184) begin
      banks_0_read_cmd_valid = 1'b1;
    end
    if(when_DataCache_l1337) begin
      banks_0_read_cmd_valid = (! (load_pipeline_stages_0_valid && (! load_pipeline_stages_0_ready)));
    end
  end

  always @(*) begin
    banks_0_read_cmd_payload = 9'bxxxxxxxxx;
    if(when_DataCache_l1184) begin
      banks_0_read_cmd_payload = {writeback_read_address[11 : 6],writeback_read_wordIndex};
    end
    if(when_DataCache_l1337) begin
      banks_0_read_cmd_payload = load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION[11 : 3];
    end
  end

  always @(*) begin
    banks_1_read_usedByWriteBack = 1'b0;
    if(when_DataCache_l1184_1) begin
      banks_1_read_usedByWriteBack = 1'b1;
    end
  end

  assign banks_1_read_rsp = _zz_banks_1_read_rsp;
  always @(*) begin
    banks_1_read_cmd_valid = 1'b0;
    if(when_DataCache_l1184_1) begin
      banks_1_read_cmd_valid = 1'b1;
    end
    if(when_DataCache_l1337_1) begin
      banks_1_read_cmd_valid = (! (load_pipeline_stages_0_valid && (! load_pipeline_stages_0_ready)));
    end
  end

  always @(*) begin
    banks_1_read_cmd_payload = 9'bxxxxxxxxx;
    if(when_DataCache_l1184_1) begin
      banks_1_read_cmd_payload = {writeback_read_address[11 : 6],writeback_read_wordIndex};
    end
    if(when_DataCache_l1337_1) begin
      banks_1_read_cmd_payload = load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION[11 : 3];
    end
  end

  always @(*) begin
    banks_2_read_usedByWriteBack = 1'b0;
    if(when_DataCache_l1184_2) begin
      banks_2_read_usedByWriteBack = 1'b1;
    end
  end

  assign banks_2_read_rsp = _zz_banks_2_read_rsp;
  always @(*) begin
    banks_2_read_cmd_valid = 1'b0;
    if(when_DataCache_l1184_2) begin
      banks_2_read_cmd_valid = 1'b1;
    end
    if(when_DataCache_l1337_2) begin
      banks_2_read_cmd_valid = (! (load_pipeline_stages_0_valid && (! load_pipeline_stages_0_ready)));
    end
  end

  always @(*) begin
    banks_2_read_cmd_payload = 9'bxxxxxxxxx;
    if(when_DataCache_l1184_2) begin
      banks_2_read_cmd_payload = {writeback_read_address[11 : 6],writeback_read_wordIndex};
    end
    if(when_DataCache_l1337_2) begin
      banks_2_read_cmd_payload = load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION[11 : 3];
    end
  end

  always @(*) begin
    banks_3_read_usedByWriteBack = 1'b0;
    if(when_DataCache_l1184_3) begin
      banks_3_read_usedByWriteBack = 1'b1;
    end
  end

  assign banks_3_read_rsp = _zz_banks_3_read_rsp;
  always @(*) begin
    banks_3_read_cmd_valid = 1'b0;
    if(when_DataCache_l1184_3) begin
      banks_3_read_cmd_valid = 1'b1;
    end
    if(when_DataCache_l1337_3) begin
      banks_3_read_cmd_valid = (! (load_pipeline_stages_0_valid && (! load_pipeline_stages_0_ready)));
    end
  end

  always @(*) begin
    banks_3_read_cmd_payload = 9'bxxxxxxxxx;
    if(when_DataCache_l1184_3) begin
      banks_3_read_cmd_payload = {writeback_read_address[11 : 6],writeback_read_wordIndex};
    end
    if(when_DataCache_l1337_3) begin
      banks_3_read_cmd_payload = load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION[11 : 3];
    end
  end

  always @(*) begin
    waysWrite_mask = 4'b0000;
    if(when_DataCache_l887) begin
      waysWrite_mask = 4'b1111;
    end
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1036) begin
        waysWrite_mask[refill_read_way] = 1'b1;
      end
    end
    if(load_ctrl_startRefill) begin
      waysWrite_mask[load_ctrl_refillWay] = 1'b1;
    end
    if(when_DataCache_l1750) begin
      waysWrite_mask[store_ctrl_refillWay] = 1'b1;
    end
    if(store_ctrl_startFlush) begin
      if(store_pipeline_stages_2_FLUSH_FREE) begin
        if(_zz_34) begin
          waysWrite_mask[0] = 1'b1;
        end
        if(_zz_store_ctrl_needFlushSel) begin
          waysWrite_mask[1] = 1'b1;
        end
        if(_zz_store_ctrl_needFlushSel_1) begin
          waysWrite_mask[2] = 1'b1;
        end
        if(_zz_store_ctrl_needFlushSel_2) begin
          waysWrite_mask[3] = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    waysWrite_address = 6'bxxxxxx;
    if(when_DataCache_l887) begin
      waysWrite_address = invalidate_counter[5:0];
    end
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1036) begin
        waysWrite_address = refill_read_rspAddress[11 : 6];
      end
    end
    if(load_ctrl_startRefill) begin
      waysWrite_address = load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[11 : 6];
    end
    if(when_DataCache_l1750) begin
      waysWrite_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 6];
    end
    if(store_ctrl_startFlush) begin
      waysWrite_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 6];
    end
  end

  always @(*) begin
    waysWrite_tag_loaded = 1'bx;
    if(when_DataCache_l887) begin
      waysWrite_tag_loaded = 1'b0;
    end
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1036) begin
        waysWrite_tag_loaded = 1'b1;
      end
    end
    if(load_ctrl_startRefill) begin
      waysWrite_tag_loaded = 1'b0;
    end
    if(when_DataCache_l1750) begin
      waysWrite_tag_loaded = 1'b0;
    end
    if(store_ctrl_startFlush) begin
      waysWrite_tag_loaded = 1'b0;
    end
  end

  always @(*) begin
    waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1036) begin
        waysWrite_tag_address = refill_read_rspAddress[31 : 12];
      end
    end
  end

  always @(*) begin
    waysWrite_tag_fault = 1'bx;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1036) begin
        waysWrite_tag_fault = refill_read_faulty;
      end
    end
  end

  assign _zz_ways_0_loadRead_rsp_loaded = _zz_ways_0_mem_port1;
  assign ways_0_loadRead_rsp_loaded = _zz_ways_0_loadRead_rsp_loaded[0];
  assign ways_0_loadRead_rsp_address = _zz_ways_0_loadRead_rsp_loaded[20 : 1];
  assign ways_0_loadRead_rsp_fault = _zz_ways_0_loadRead_rsp_loaded[21];
  assign _zz_ways_0_storeRead_rsp_loaded = _zz_ways_0_mem_port2;
  assign ways_0_storeRead_rsp_loaded = _zz_ways_0_storeRead_rsp_loaded[0];
  assign ways_0_storeRead_rsp_address = _zz_ways_0_storeRead_rsp_loaded[20 : 1];
  assign ways_0_storeRead_rsp_fault = _zz_ways_0_storeRead_rsp_loaded[21];
  assign _zz_ways_1_loadRead_rsp_loaded = _zz_ways_1_mem_port1;
  assign ways_1_loadRead_rsp_loaded = _zz_ways_1_loadRead_rsp_loaded[0];
  assign ways_1_loadRead_rsp_address = _zz_ways_1_loadRead_rsp_loaded[20 : 1];
  assign ways_1_loadRead_rsp_fault = _zz_ways_1_loadRead_rsp_loaded[21];
  assign _zz_ways_1_storeRead_rsp_loaded = _zz_ways_1_mem_port2;
  assign ways_1_storeRead_rsp_loaded = _zz_ways_1_storeRead_rsp_loaded[0];
  assign ways_1_storeRead_rsp_address = _zz_ways_1_storeRead_rsp_loaded[20 : 1];
  assign ways_1_storeRead_rsp_fault = _zz_ways_1_storeRead_rsp_loaded[21];
  assign _zz_ways_2_loadRead_rsp_loaded = _zz_ways_2_mem_port1;
  assign ways_2_loadRead_rsp_loaded = _zz_ways_2_loadRead_rsp_loaded[0];
  assign ways_2_loadRead_rsp_address = _zz_ways_2_loadRead_rsp_loaded[20 : 1];
  assign ways_2_loadRead_rsp_fault = _zz_ways_2_loadRead_rsp_loaded[21];
  assign _zz_ways_2_storeRead_rsp_loaded = _zz_ways_2_mem_port2;
  assign ways_2_storeRead_rsp_loaded = _zz_ways_2_storeRead_rsp_loaded[0];
  assign ways_2_storeRead_rsp_address = _zz_ways_2_storeRead_rsp_loaded[20 : 1];
  assign ways_2_storeRead_rsp_fault = _zz_ways_2_storeRead_rsp_loaded[21];
  assign _zz_ways_3_loadRead_rsp_loaded = _zz_ways_3_mem_port1;
  assign ways_3_loadRead_rsp_loaded = _zz_ways_3_loadRead_rsp_loaded[0];
  assign ways_3_loadRead_rsp_address = _zz_ways_3_loadRead_rsp_loaded[20 : 1];
  assign ways_3_loadRead_rsp_fault = _zz_ways_3_loadRead_rsp_loaded[21];
  assign _zz_ways_3_storeRead_rsp_loaded = _zz_ways_3_mem_port2;
  assign ways_3_storeRead_rsp_loaded = _zz_ways_3_storeRead_rsp_loaded[0];
  assign ways_3_storeRead_rsp_address = _zz_ways_3_storeRead_rsp_loaded[20 : 1];
  assign ways_3_storeRead_rsp_fault = _zz_ways_3_storeRead_rsp_loaded[21];
  always @(*) begin
    status_write_valid = 1'b0;
    if(load_ctrl_startRefill) begin
      status_write_valid = 1'b1;
    end
    if(when_DataCache_l1725) begin
      status_write_valid = 1'b1;
    end
  end

  always @(*) begin
    status_write_payload_address = 6'bxxxxxx;
    if(load_ctrl_startRefill) begin
      status_write_payload_address = load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[11 : 6];
    end
    if(when_DataCache_l1725) begin
      status_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 6];
    end
  end

  always @(*) begin
    status_write_payload_data_0_dirty = 1'bx;
    if(load_ctrl_startRefill) begin
      status_write_payload_data_0_dirty = load_pipeline_stages_2_STATUS_0_dirty;
      if(_zz_32[0]) begin
        status_write_payload_data_0_dirty = 1'b0;
      end
    end
    if(when_DataCache_l1725) begin
      status_write_payload_data_0_dirty = store_pipeline_stages_2_STATUS_0_dirty;
    end
    if(when_DataCache_l1750) begin
      case(store_ctrl_refillWay)
        2'b00 : begin
          status_write_payload_data_0_dirty = 1'b0;
        end
        2'b01 : begin
        end
        2'b10 : begin
        end
        default : begin
        end
      endcase
    end
    if(store_ctrl_setDirty) begin
      if(store_pipeline_stages_2_WAYS_HITS[0]) begin
        status_write_payload_data_0_dirty = 1'b1;
      end
    end
    if(store_ctrl_startFlush) begin
      if(_zz_34) begin
        status_write_payload_data_0_dirty = 1'b0;
      end
    end
  end

  always @(*) begin
    status_write_payload_data_1_dirty = 1'bx;
    if(load_ctrl_startRefill) begin
      status_write_payload_data_1_dirty = load_pipeline_stages_2_STATUS_1_dirty;
      if(_zz_32[1]) begin
        status_write_payload_data_1_dirty = 1'b0;
      end
    end
    if(when_DataCache_l1725) begin
      status_write_payload_data_1_dirty = store_pipeline_stages_2_STATUS_1_dirty;
    end
    if(when_DataCache_l1750) begin
      case(store_ctrl_refillWay)
        2'b00 : begin
        end
        2'b01 : begin
          status_write_payload_data_1_dirty = 1'b0;
        end
        2'b10 : begin
        end
        default : begin
        end
      endcase
    end
    if(store_ctrl_setDirty) begin
      if(_zz_store_ctrl_wayId) begin
        status_write_payload_data_1_dirty = 1'b1;
      end
    end
    if(store_ctrl_startFlush) begin
      if(_zz_store_ctrl_needFlushSel) begin
        status_write_payload_data_1_dirty = 1'b0;
      end
    end
  end

  always @(*) begin
    status_write_payload_data_2_dirty = 1'bx;
    if(load_ctrl_startRefill) begin
      status_write_payload_data_2_dirty = load_pipeline_stages_2_STATUS_2_dirty;
      if(_zz_32[2]) begin
        status_write_payload_data_2_dirty = 1'b0;
      end
    end
    if(when_DataCache_l1725) begin
      status_write_payload_data_2_dirty = store_pipeline_stages_2_STATUS_2_dirty;
    end
    if(when_DataCache_l1750) begin
      case(store_ctrl_refillWay)
        2'b00 : begin
        end
        2'b01 : begin
        end
        2'b10 : begin
          status_write_payload_data_2_dirty = 1'b0;
        end
        default : begin
        end
      endcase
    end
    if(store_ctrl_setDirty) begin
      if(_zz_store_ctrl_wayId_1) begin
        status_write_payload_data_2_dirty = 1'b1;
      end
    end
    if(store_ctrl_startFlush) begin
      if(_zz_store_ctrl_needFlushSel_1) begin
        status_write_payload_data_2_dirty = 1'b0;
      end
    end
  end

  always @(*) begin
    status_write_payload_data_3_dirty = 1'bx;
    if(load_ctrl_startRefill) begin
      status_write_payload_data_3_dirty = load_pipeline_stages_2_STATUS_3_dirty;
      if(_zz_32[3]) begin
        status_write_payload_data_3_dirty = 1'b0;
      end
    end
    if(when_DataCache_l1725) begin
      status_write_payload_data_3_dirty = store_pipeline_stages_2_STATUS_3_dirty;
    end
    if(when_DataCache_l1750) begin
      case(store_ctrl_refillWay)
        2'b00 : begin
        end
        2'b01 : begin
        end
        2'b10 : begin
        end
        default : begin
          status_write_payload_data_3_dirty = 1'b0;
        end
      endcase
    end
    if(store_ctrl_setDirty) begin
      if(_zz_store_ctrl_wayId_2) begin
        status_write_payload_data_3_dirty = 1'b1;
      end
    end
    if(store_ctrl_startFlush) begin
      if(_zz_store_ctrl_needFlushSel_2) begin
        status_write_payload_data_3_dirty = 1'b0;
      end
    end
  end

  assign _zz_status_loadRead_rsp_0_dirty = _zz_status_mem_port1;
  assign status_loadRead_rsp_0_dirty = _zz_status_loadRead_rsp_0_dirty_1[0];
  assign status_loadRead_rsp_1_dirty = _zz_status_loadRead_rsp_1_dirty[0];
  assign status_loadRead_rsp_2_dirty = _zz_status_loadRead_rsp_2_dirty[0];
  assign status_loadRead_rsp_3_dirty = _zz_status_loadRead_rsp_3_dirty[0];
  assign _zz_status_storeRead_rsp_0_dirty = _zz_status_mem_port2;
  assign status_storeRead_rsp_0_dirty = _zz_status_storeRead_rsp_0_dirty_1[0];
  assign status_storeRead_rsp_1_dirty = _zz_status_storeRead_rsp_1_dirty[0];
  assign status_storeRead_rsp_2_dirty = _zz_status_storeRead_rsp_2_dirty[0];
  assign status_storeRead_rsp_3_dirty = _zz_status_storeRead_rsp_3_dirty[0];
  assign wayRandom_willClear = 1'b0;
  assign wayRandom_willOverflowIfInc = (wayRandom_value == 2'b11);
  assign wayRandom_willOverflow = (wayRandom_willOverflowIfInc && wayRandom_willIncrement);
  always @(*) begin
    wayRandom_valueNext = (wayRandom_value + _zz_wayRandom_valueNext);
    if(wayRandom_willClear) begin
      wayRandom_valueNext = 2'b00;
    end
  end

  assign wayRandom_willIncrement = 1'b1;
  always @(*) begin
    plru_write_valid = (plru_fromLoad_valid || plru_fromStore_valid);
    if(when_DataCache_l896) begin
      plru_write_valid = 1'b1;
    end
  end

  always @(*) begin
    plru_write_payload_address = (plru_fromLoad_valid ? plru_fromLoad_payload_address : plru_fromStore_payload_address);
    if(when_DataCache_l896) begin
      plru_write_payload_address = invalidate_counter[5:0];
    end
  end

  always @(*) begin
    plru_write_payload_data_0 = (plru_fromLoad_valid ? plru_fromLoad_payload_data_0 : plru_fromStore_payload_data_0);
    if(when_DataCache_l896) begin
      plru_write_payload_data_0 = _zz_plru_write_payload_data_0[0 : 0];
    end
  end

  always @(*) begin
    plru_write_payload_data_1 = (plru_fromLoad_valid ? plru_fromLoad_payload_data_1 : plru_fromStore_payload_data_1);
    if(when_DataCache_l896) begin
      plru_write_payload_data_1 = _zz_plru_write_payload_data_0[2 : 1];
    end
  end

  assign invalidate_done = invalidate_counter[6];
  always @(*) begin
    invalidate_reservation_take = 1'b0;
    if(when_DataCache_l887) begin
      invalidate_reservation_take = 1'b1;
    end
  end

  assign when_DataCache_l887 = ((! invalidate_done) && invalidate_reservation_win);
  assign when_DataCache_l896 = ((! invalidate_done) && invalidate_firstEver);
  assign _zz_plru_write_payload_data_0 = 3'b000;
  assign refill_slots_0_loadedDone = (refill_slots_0_loadedCounter == 1'b1);
  assign when_DataCache_l933 = (refill_slots_0_loadedDone && 1'b1);
  assign refill_slots_0_free = (! refill_slots_0_valid);
  assign refill_slots_1_loadedDone = (refill_slots_1_loadedCounter == 1'b1);
  assign when_DataCache_l933_1 = (refill_slots_1_loadedDone && 1'b1);
  assign refill_slots_1_free = (! refill_slots_1_valid);
  assign _zz_refill_free = {refill_slots_1_free,refill_slots_0_free};
  assign refill_free = {_zz_refill_free_1[1],refill_slots_0_free};
  assign refill_full = ((! refill_slots_0_free) && (! refill_slots_1_free));
  always @(*) begin
    refill_push_valid = 1'b0;
    if(when_DataCache_l1471) begin
      refill_push_valid = 1'b1;
    end
    if(when_DataCache_l1750) begin
      refill_push_valid = 1'b1;
    end
  end

  always @(*) begin
    refill_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_DataCache_l1471) begin
      refill_push_payload_address = load_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
    end
    if(when_DataCache_l1750) begin
      refill_push_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
    end
  end

  always @(*) begin
    refill_push_payload_way = 2'bxx;
    if(load_ctrl_askUpgrade) begin
      refill_push_payload_way = load_ctrl_wayId;
    end else begin
      refill_push_payload_way = load_ctrl_refillWay;
    end
    if(when_DataCache_l1750) begin
      refill_push_payload_way = store_ctrl_refillWay;
    end
  end

  always @(*) begin
    refill_push_payload_victim = 2'bxx;
    if(load_ctrl_askUpgrade) begin
      refill_push_payload_victim = 2'b00;
    end else begin
      refill_push_payload_victim = ((load_ctrl_refillWayNeedWriteback && _zz_refill_push_payload_victim) ? writeback_free : 2'b00);
    end
    if(when_DataCache_l1750) begin
      refill_push_payload_victim = (((store_ctrl_replacedWayNeedWriteback && store_ctrl_askRefill) && _zz_refill_push_payload_victim_1) ? writeback_free : 2'b00);
    end
  end

  always @(*) begin
    refill_push_payload_unique = 1'bx;
    if(when_DataCache_l1471) begin
      refill_push_payload_unique = load_pipeline_stages_2_NEED_UNIQUE;
    end
    if(when_DataCache_l1750) begin
      refill_push_payload_unique = 1'b1;
    end
  end

  always @(*) begin
    refill_push_payload_data = 1'bx;
    if(when_DataCache_l1471) begin
      refill_push_payload_data = load_ctrl_askRefill;
    end
    if(when_DataCache_l1750) begin
      refill_push_payload_data = store_ctrl_askRefill;
    end
  end

  assign when_DataCache_l960 = refill_free[0];
  assign _zz_27 = refill_free[0];
  assign _zz_28 = refill_free[1];
  assign when_DataCache_l960_1 = refill_free[1];
  assign refill_read_arbiter_slotsWithId_0_0 = (((refill_slots_0_valid && (! refill_slots_0_cmdSent)) && (refill_slots_0_victim == 2'b00)) && (refill_slots_0_writebackHazards == 2'b00));
  assign refill_read_arbiter_slotsWithId_1_0 = (((refill_slots_1_valid && (! refill_slots_1_cmdSent)) && (refill_slots_1_victim == 2'b00)) && (refill_slots_1_writebackHazards == 2'b00));
  assign refill_read_arbiter_hits = {refill_read_arbiter_slotsWithId_1_0,refill_read_arbiter_slotsWithId_0_0};
  assign refill_read_arbiter_hit = (|refill_read_arbiter_hits);
  always @(*) begin
    refill_read_arbiter_oh = (refill_read_arbiter_hits & {((refill_read_arbiter_hits[0] & refill_slots_1_priority) == 1'b0),((refill_read_arbiter_hits[1] & refill_slots_0_priority) == 1'b0)});
    if(when_DataCache_l910) begin
      refill_read_arbiter_oh = refill_read_arbiter_lock;
    end
  end

  assign _zz_refill_read_arbiter_sel = refill_read_arbiter_oh[1];
  assign refill_read_arbiter_sel = _zz_refill_read_arbiter_sel;
  assign when_DataCache_l910 = (|refill_read_arbiter_lock);
  assign refill_read_writebackHazard = (|refill_read_writebackHazards);
  assign io_mem_read_cmd_fire = (io_mem_read_cmd_valid && io_mem_read_cmd_ready);
  assign when_DataCache_l985 = (io_mem_read_cmd_fire || refill_read_writebackHazard);
  assign refill_read_cmdAddress = {_zz_refill_read_cmdAddress,6'h00};
  assign io_mem_read_cmd_valid = (refill_read_arbiter_hit && (! refill_read_writebackHazard));
  assign io_mem_read_cmd_payload_id = refill_read_arbiter_sel;
  assign io_mem_read_cmd_payload_address = refill_read_cmdAddress;
  assign when_DataCache_l997 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign when_DataCache_l997_1 = (io_mem_read_cmd_ready && (! refill_read_writebackHazard));
  assign refill_read_rspAddress = _zz_refill_read_rspAddress;
  assign refill_read_way = _zz_refill_read_way;
  assign refill_read_rspWithData = 1'b1;
  always @(*) begin
    refill_read_bankWriteNotif = 4'b0000;
    refill_read_bankWriteNotif[0] = ((io_mem_read_rsp_valid && refill_read_rspWithData) && (refill_read_way == 2'b00));
    refill_read_bankWriteNotif[1] = ((io_mem_read_rsp_valid && refill_read_rspWithData) && (refill_read_way == 2'b01));
    refill_read_bankWriteNotif[2] = ((io_mem_read_rsp_valid && refill_read_rspWithData) && (refill_read_way == 2'b10));
    refill_read_bankWriteNotif[3] = ((io_mem_read_rsp_valid && refill_read_rspWithData) && (refill_read_way == 2'b11));
  end

  always @(*) begin
    banks_0_write_valid = refill_read_bankWriteNotif[0];
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774) begin
        banks_0_write_valid = (2'b00 == store_ctrl_wayId);
      end
    end
  end

  always @(*) begin
    banks_0_write_payload_address = {refill_read_rspAddress[11 : 6],refill_read_wordIndex};
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774) begin
        banks_0_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 3];
      end
    end
  end

  always @(*) begin
    banks_0_write_payload_data = io_mem_read_rsp_payload_data;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774) begin
        banks_0_write_payload_data[31 : 0] = store_pipeline_stages_2_CPU_WORD;
        banks_0_write_payload_data[63 : 32] = store_pipeline_stages_2_CPU_WORD;
      end
    end
  end

  always @(*) begin
    banks_0_write_payload_mask = 8'hff;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774) begin
        banks_0_write_payload_mask = 8'h00;
        if(_zz_35[0]) begin
          banks_0_write_payload_mask[3 : 0] = store_pipeline_stages_2_CPU_MASK;
        end
        if(_zz_35[1]) begin
          banks_0_write_payload_mask[7 : 4] = store_pipeline_stages_2_CPU_MASK;
        end
      end
    end
  end

  always @(*) begin
    banks_1_write_valid = refill_read_bankWriteNotif[1];
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_1) begin
        banks_1_write_valid = (2'b01 == store_ctrl_wayId);
      end
    end
  end

  always @(*) begin
    banks_1_write_payload_address = {refill_read_rspAddress[11 : 6],refill_read_wordIndex};
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_1) begin
        banks_1_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 3];
      end
    end
  end

  always @(*) begin
    banks_1_write_payload_data = io_mem_read_rsp_payload_data;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_1) begin
        banks_1_write_payload_data[31 : 0] = store_pipeline_stages_2_CPU_WORD;
        banks_1_write_payload_data[63 : 32] = store_pipeline_stages_2_CPU_WORD;
      end
    end
  end

  always @(*) begin
    banks_1_write_payload_mask = 8'hff;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_1) begin
        banks_1_write_payload_mask = 8'h00;
        if(_zz_36[0]) begin
          banks_1_write_payload_mask[3 : 0] = store_pipeline_stages_2_CPU_MASK;
        end
        if(_zz_36[1]) begin
          banks_1_write_payload_mask[7 : 4] = store_pipeline_stages_2_CPU_MASK;
        end
      end
    end
  end

  always @(*) begin
    banks_2_write_valid = refill_read_bankWriteNotif[2];
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_2) begin
        banks_2_write_valid = (2'b10 == store_ctrl_wayId);
      end
    end
  end

  always @(*) begin
    banks_2_write_payload_address = {refill_read_rspAddress[11 : 6],refill_read_wordIndex};
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_2) begin
        banks_2_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 3];
      end
    end
  end

  always @(*) begin
    banks_2_write_payload_data = io_mem_read_rsp_payload_data;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_2) begin
        banks_2_write_payload_data[31 : 0] = store_pipeline_stages_2_CPU_WORD;
        banks_2_write_payload_data[63 : 32] = store_pipeline_stages_2_CPU_WORD;
      end
    end
  end

  always @(*) begin
    banks_2_write_payload_mask = 8'hff;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_2) begin
        banks_2_write_payload_mask = 8'h00;
        if(_zz_37[0]) begin
          banks_2_write_payload_mask[3 : 0] = store_pipeline_stages_2_CPU_MASK;
        end
        if(_zz_37[1]) begin
          banks_2_write_payload_mask[7 : 4] = store_pipeline_stages_2_CPU_MASK;
        end
      end
    end
  end

  always @(*) begin
    banks_3_write_valid = refill_read_bankWriteNotif[3];
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_3) begin
        banks_3_write_valid = (2'b11 == store_ctrl_wayId);
      end
    end
  end

  always @(*) begin
    banks_3_write_payload_address = {refill_read_rspAddress[11 : 6],refill_read_wordIndex};
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_3) begin
        banks_3_write_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 3];
      end
    end
  end

  always @(*) begin
    banks_3_write_payload_data = io_mem_read_rsp_payload_data;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_3) begin
        banks_3_write_payload_data[31 : 0] = store_pipeline_stages_2_CPU_WORD;
        banks_3_write_payload_data[63 : 32] = store_pipeline_stages_2_CPU_WORD;
      end
    end
  end

  always @(*) begin
    banks_3_write_payload_mask = 8'hff;
    if(store_ctrl_writeCache) begin
      if(when_DataCache_l1774_3) begin
        banks_3_write_payload_mask = 8'h00;
        if(_zz_38[0]) begin
          banks_3_write_payload_mask[3 : 0] = store_pipeline_stages_2_CPU_MASK;
        end
        if(_zz_38[1]) begin
          banks_3_write_payload_mask[7 : 4] = store_pipeline_stages_2_CPU_MASK;
        end
      end
    end
  end

  assign when_DataCache_l1025 = (io_mem_read_rsp_valid && io_mem_read_rsp_payload_error);
  always @(*) begin
    refill_read_fire = 1'b0;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1036) begin
        refill_read_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    refill_read_reservation_take = 1'b0;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1036) begin
        refill_read_reservation_take = 1'b1;
      end
    end
  end

  assign refill_read_faulty = (refill_read_hadError || io_mem_read_rsp_payload_error);
  always @(*) begin
    io_refillCompletions = 2'b00;
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1036) begin
        io_refillCompletions[io_mem_read_rsp_payload_id] = 1'b1;
      end
    end
  end

  assign io_mem_read_rsp_ready = 1'b1;
  assign when_DataCache_l1036 = ((refill_read_wordIndex == 3'b111) || (! refill_read_rspWithData));
  always @(*) begin
    writeback_slots_0_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        1'b0 : begin
          writeback_slots_0_fire = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  assign writeback_slots_0_free = (! writeback_slots_0_valid);
  always @(*) begin
    refill_read_writebackHazards[0] = (writeback_slots_0_valid && (writeback_slots_0_address[31 : 6] == refill_read_cmdAddress[31 : 6]));
    refill_read_writebackHazards[1] = (writeback_slots_1_valid && (writeback_slots_1_address[31 : 6] == refill_read_cmdAddress[31 : 6]));
  end

  always @(*) begin
    writeback_slots_1_fire = 1'b0;
    if(io_mem_write_rsp_valid) begin
      case(io_mem_write_rsp_payload_id)
        1'b0 : begin
        end
        default : begin
          writeback_slots_1_fire = 1'b1;
        end
      endcase
    end
  end

  assign writeback_slots_1_free = (! writeback_slots_1_valid);
  assign io_writebackBusy = ({writeback_slots_1_valid,writeback_slots_0_valid} != 2'b00);
  assign _zz_writeback_free = {writeback_slots_1_free,writeback_slots_0_free};
  assign writeback_free = {_zz_writeback_free_1[1],writeback_slots_0_free};
  assign writeback_full = ((! writeback_slots_0_free) && (! writeback_slots_1_free));
  always @(*) begin
    writeback_push_valid = 1'b0;
    if(load_ctrl_startRefill) begin
      writeback_push_valid = load_ctrl_refillWayNeedWriteback;
    end
    if(when_DataCache_l1732) begin
      writeback_push_valid = (store_ctrl_replacedWayNeedWriteback || store_ctrl_startFlush);
    end
  end

  always @(*) begin
    writeback_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(load_ctrl_startRefill) begin
      writeback_push_payload_address = ({6'd0,{_zz_writeback_push_payload_address,load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[11 : 6]}} <<< 3'd6);
    end
    if(when_DataCache_l1732) begin
      writeback_push_payload_address = ({6'd0,{_zz_writeback_push_payload_address_1,store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 6]}} <<< 3'd6);
    end
  end

  always @(*) begin
    writeback_push_payload_way = 2'bxx;
    if(load_ctrl_startRefill) begin
      writeback_push_payload_way = load_ctrl_refillWay;
    end
    if(when_DataCache_l1732) begin
      writeback_push_payload_way = (store_pipeline_stages_2_FLUSH ? store_ctrl_needFlushSel : store_ctrl_refillWay);
    end
  end

  assign when_DataCache_l1127 = writeback_free[0];
  assign when_DataCache_l1127_1 = writeback_free[1];
  assign writeback_read_arbiter_slotsWithId_0_0 = (writeback_slots_0_valid && (! writeback_slots_0_readCmdDone));
  assign writeback_read_arbiter_slotsWithId_1_0 = (writeback_slots_1_valid && (! writeback_slots_1_readCmdDone));
  assign writeback_read_arbiter_hits = {writeback_read_arbiter_slotsWithId_1_0,writeback_read_arbiter_slotsWithId_0_0};
  assign writeback_read_arbiter_hit = (|writeback_read_arbiter_hits);
  always @(*) begin
    writeback_read_arbiter_oh = (writeback_read_arbiter_hits & {((writeback_read_arbiter_hits[0] & writeback_slots_1_priority) == 1'b0),((writeback_read_arbiter_hits[1] & writeback_slots_0_priority) == 1'b0)});
    if(when_DataCache_l910_1) begin
      writeback_read_arbiter_oh = writeback_read_arbiter_lock;
    end
  end

  assign _zz_writeback_read_arbiter_sel = writeback_read_arbiter_oh[1];
  assign writeback_read_arbiter_sel = _zz_writeback_read_arbiter_sel;
  assign when_DataCache_l910_1 = (|writeback_read_arbiter_lock);
  assign writeback_read_address = _zz_writeback_read_address;
  assign writeback_read_way = _zz_writeback_read_way;
  assign writeback_read_slotRead_valid = writeback_read_arbiter_hit;
  assign writeback_read_slotRead_payload_id = writeback_read_arbiter_sel;
  assign writeback_read_slotRead_payload_wordIndex = writeback_read_wordIndex;
  assign writeback_read_slotRead_payload_way = writeback_read_way;
  assign writeback_read_slotRead_payload_last = (writeback_read_wordIndex == 3'b111);
  assign when_DataCache_l1174 = (writeback_read_slotRead_valid && writeback_read_slotRead_payload_last);
  assign when_DataCache_l1184 = (writeback_read_slotRead_valid && (writeback_read_way == 2'b00));
  assign when_DataCache_l1184_1 = (writeback_read_slotRead_valid && (writeback_read_way == 2'b01));
  assign when_DataCache_l1184_2 = (writeback_read_slotRead_valid && (writeback_read_way == 2'b10));
  assign when_DataCache_l1184_3 = (writeback_read_slotRead_valid && (writeback_read_way == 2'b11));
  assign writeback_read_readedData = _zz_writeback_read_readedData;
  assign _zz_when_MultiportRam_l328_1 = {writeback_read_slotReadLast_payload_id,writeback_read_slotReadLast_payload_wordIndex};
  assign writeback_write_arbiter_slotsWithId_0_0 = ((writeback_slots_0_valid && writeback_slots_0_victimBufferReady) && (! writeback_slots_0_writeCmdDone));
  assign writeback_write_arbiter_slotsWithId_1_0 = ((writeback_slots_1_valid && writeback_slots_1_victimBufferReady) && (! writeback_slots_1_writeCmdDone));
  assign writeback_write_arbiter_hits = {writeback_write_arbiter_slotsWithId_1_0,writeback_write_arbiter_slotsWithId_0_0};
  assign writeback_write_arbiter_hit = (|writeback_write_arbiter_hits);
  always @(*) begin
    writeback_write_arbiter_oh = (writeback_write_arbiter_hits & {((writeback_write_arbiter_hits[0] & writeback_slots_1_priority) == 1'b0),((writeback_write_arbiter_hits[1] & writeback_slots_0_priority) == 1'b0)});
    if(when_DataCache_l910_2) begin
      writeback_write_arbiter_oh = writeback_write_arbiter_lock;
    end
  end

  assign _zz_writeback_write_arbiter_sel = writeback_write_arbiter_oh[1];
  assign writeback_write_arbiter_sel = _zz_writeback_write_arbiter_sel;
  assign when_DataCache_l910_2 = (|writeback_write_arbiter_lock);
  assign writeback_write_last = (writeback_write_wordIndex == 3'b111);
  assign writeback_write_bufferRead_valid = writeback_write_arbiter_hit;
  assign writeback_write_bufferRead_payload_id = writeback_write_arbiter_sel;
  assign writeback_write_bufferRead_payload_last = writeback_write_last;
  assign writeback_write_bufferRead_payload_address = _zz_writeback_write_bufferRead_payload_address;
  assign writeback_write_bufferRead_fire = (writeback_write_bufferRead_valid && writeback_write_bufferRead_ready);
  assign when_DataCache_l1252 = (writeback_write_bufferRead_fire && writeback_write_last);
  always @(*) begin
    writeback_write_bufferRead_ready = writeback_write_cmd_ready;
    if(when_Stream_l369) begin
      writeback_write_bufferRead_ready = 1'b1;
    end
  end

  assign when_Stream_l369 = (! writeback_write_cmd_valid);
  assign writeback_write_cmd_valid = writeback_write_bufferRead_rValid;
  assign writeback_write_cmd_payload_id = writeback_write_bufferRead_rData_id;
  assign writeback_write_cmd_payload_address = writeback_write_bufferRead_rData_address;
  assign writeback_write_cmd_payload_last = writeback_write_bufferRead_rData_last;
  assign _zz_when_MultiportRam_l328_2 = {writeback_write_bufferRead_payload_id,writeback_write_wordIndex};
  assign writeback_write_word = _zz_writeback_write_word;
  assign io_mem_write_cmd_valid = writeback_write_cmd_valid;
  assign writeback_write_cmd_ready = io_mem_write_cmd_ready;
  assign io_mem_write_cmd_payload_fragment_address = writeback_write_cmd_payload_address;
  assign io_mem_write_cmd_payload_fragment_data = writeback_write_word;
  assign io_mem_write_cmd_payload_fragment_id = writeback_write_cmd_payload_id;
  assign io_mem_write_cmd_payload_last = writeback_write_cmd_payload_last;
  assign _zz_load_pipeline_stages_0_throwRequest_DataCache_l1301 = io_load_cancels[0];
  assign load_pipeline_stages_0_throwRequest_DataCache_l1301 = _zz_load_pipeline_stages_0_throwRequest_DataCache_l1301;
  assign _zz_load_pipeline_stages_1_throwRequest_DataCache_l1301 = io_load_cancels[1];
  assign load_pipeline_stages_1_throwRequest_DataCache_l1301 = _zz_load_pipeline_stages_1_throwRequest_DataCache_l1301;
  assign load_pipeline_stages_2_throwRequest_DataCache_l1301 = io_load_cancels[2];
  assign load_pipeline_stages_1_WAYS_HAZARD_overloaded = (load_pipeline_stages_1_WAYS_HAZARD | ((waysWrite_addressLast == load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[11 : 6]) ? waysWrite_maskLast : 4'b0000));
  assign load_pipeline_stages_2_WAYS_HAZARD_overloaded = (load_pipeline_stages_2_WAYS_HAZARD | ((waysWrite_addressLast == load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[11 : 6]) ? waysWrite_maskLast : 4'b0000));
  assign io_load_cmd_ready = 1'b1;
  assign load_pipeline_stages_0_valid = io_load_cmd_valid;
  assign load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION = io_load_cmd_payload_virtual;
  assign load_pipeline_stages_0_REDO_ON_DATA_HAZARD = io_load_cmd_payload_redoOnDataHazard;
  assign load_pipeline_stages_0_WAYS_HAZARD = 4'b0000;
  assign load_pipeline_stages_0_UNLOCKED = io_load_cmd_payload_unlocked;
  assign load_pipeline_stages_0_NEED_UNIQUE = io_load_cmd_payload_unique;
  always @(*) begin
    load_pipeline_stages_0_BANK_BUSY[0] = banks_0_read_usedByWriteBack;
    load_pipeline_stages_0_BANK_BUSY[1] = banks_1_read_usedByWriteBack;
    load_pipeline_stages_0_BANK_BUSY[2] = banks_2_read_usedByWriteBack;
    load_pipeline_stages_0_BANK_BUSY[3] = banks_3_read_usedByWriteBack;
  end

  assign when_DataCache_l1337 = (! load_pipeline_stages_0_BANK_BUSY[0]);
  always @(*) begin
    load_pipeline_stages_0_BANK_BUSY_overloaded[0] = (load_pipeline_stages_0_BANK_BUSY[0] || (banks_0_write_valid && load_pipeline_stages_0_REDO_ON_DATA_HAZARD));
    load_pipeline_stages_0_BANK_BUSY_overloaded[1] = (load_pipeline_stages_0_BANK_BUSY[1] || (banks_1_write_valid && load_pipeline_stages_0_REDO_ON_DATA_HAZARD));
    load_pipeline_stages_0_BANK_BUSY_overloaded[2] = (load_pipeline_stages_0_BANK_BUSY[2] || (banks_2_write_valid && load_pipeline_stages_0_REDO_ON_DATA_HAZARD));
    load_pipeline_stages_0_BANK_BUSY_overloaded[3] = (load_pipeline_stages_0_BANK_BUSY[3] || (banks_3_write_valid && load_pipeline_stages_0_REDO_ON_DATA_HAZARD));
  end

  assign load_pipeline_stages_1_BANKS_WORDS_0 = banks_0_read_rsp;
  always @(*) begin
    load_pipeline_stages_1_BANK_BUSY_REMAPPED[0] = load_pipeline_stages_1_BANK_BUSY[2'b00];
    load_pipeline_stages_1_BANK_BUSY_REMAPPED[1] = load_pipeline_stages_1_BANK_BUSY[2'b01];
    load_pipeline_stages_1_BANK_BUSY_REMAPPED[2] = load_pipeline_stages_1_BANK_BUSY[2'b10];
    load_pipeline_stages_1_BANK_BUSY_REMAPPED[3] = load_pipeline_stages_1_BANK_BUSY[2'b11];
  end

  assign load_pipeline_stages_1_BANKS_MUXES_0 = _zz_load_pipeline_stages_1_BANKS_MUXES_0;
  assign when_DataCache_l1337_1 = (! load_pipeline_stages_0_BANK_BUSY[1]);
  assign load_pipeline_stages_1_BANKS_WORDS_1 = banks_1_read_rsp;
  assign load_pipeline_stages_1_BANKS_MUXES_1 = _zz_load_pipeline_stages_1_BANKS_MUXES_1;
  assign when_DataCache_l1337_2 = (! load_pipeline_stages_0_BANK_BUSY[2]);
  assign load_pipeline_stages_1_BANKS_WORDS_2 = banks_2_read_rsp;
  assign load_pipeline_stages_1_BANKS_MUXES_2 = _zz_load_pipeline_stages_1_BANKS_MUXES_2;
  assign when_DataCache_l1337_3 = (! load_pipeline_stages_0_BANK_BUSY[3]);
  assign load_pipeline_stages_1_BANKS_WORDS_3 = banks_3_read_rsp;
  assign load_pipeline_stages_1_BANKS_MUXES_3 = _zz_load_pipeline_stages_1_BANKS_MUXES_3;
  assign _zz_load_pipeline_stages_2_CPU_WORD = load_pipeline_stages_2_WAYS_HITS[1];
  assign _zz_load_pipeline_stages_2_CPU_WORD_1 = load_pipeline_stages_2_WAYS_HITS[2];
  assign _zz_load_pipeline_stages_2_CPU_WORD_2 = load_pipeline_stages_2_WAYS_HITS[3];
  assign load_pipeline_stages_2_CPU_WORD = (((load_pipeline_stages_2_WAYS_HITS[0] ? load_pipeline_stages_2_BANKS_MUXES_0 : 32'h00000000) | (_zz_load_pipeline_stages_2_CPU_WORD ? load_pipeline_stages_2_BANKS_MUXES_1 : 32'h00000000)) | ((_zz_load_pipeline_stages_2_CPU_WORD_1 ? load_pipeline_stages_2_BANKS_MUXES_2 : 32'h00000000) | (_zz_load_pipeline_stages_2_CPU_WORD_2 ? load_pipeline_stages_2_BANKS_MUXES_3 : 32'h00000000)));
  assign load_pipeline_stages_1_ADDRESS_POST_TRANSLATION = io_load_translated_physical;
  assign load_pipeline_stages_1_ABORD = io_load_translated_abord;
  assign _zz_load_pipeline_stages_1_PLRU_0 = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[11 : 6];
  assign _zz_load_pipeline_stages_1_PLRU_0_1 = _zz_plru_ram_port1;
  assign load_pipeline_stages_1_PLRU_0 = _zz_load_pipeline_stages_1_PLRU_0_1[0 : 0];
  assign load_pipeline_stages_1_PLRU_1 = _zz_load_pipeline_stages_1_PLRU_0_1[2 : 1];
  assign ways_0_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign ways_0_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[11 : 6];
  assign load_pipeline_stages_1_WAYS_TAGS_0_loaded = ways_0_loadRead_rsp_loaded;
  assign load_pipeline_stages_1_WAYS_TAGS_0_address = ways_0_loadRead_rsp_address;
  assign load_pipeline_stages_1_WAYS_TAGS_0_fault = ways_0_loadRead_rsp_fault;
  always @(*) begin
    load_pipeline_stages_1_WAYS_HITS[0] = (load_pipeline_stages_1_WAYS_TAGS_0_loaded && (load_pipeline_stages_1_WAYS_TAGS_0_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 12]));
    load_pipeline_stages_1_WAYS_HITS[1] = (load_pipeline_stages_1_WAYS_TAGS_1_loaded && (load_pipeline_stages_1_WAYS_TAGS_1_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 12]));
    load_pipeline_stages_1_WAYS_HITS[2] = (load_pipeline_stages_1_WAYS_TAGS_2_loaded && (load_pipeline_stages_1_WAYS_TAGS_2_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 12]));
    load_pipeline_stages_1_WAYS_HITS[3] = (load_pipeline_stages_1_WAYS_TAGS_3_loaded && (load_pipeline_stages_1_WAYS_TAGS_3_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 12]));
  end

  assign ways_1_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign ways_1_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[11 : 6];
  assign load_pipeline_stages_1_WAYS_TAGS_1_loaded = ways_1_loadRead_rsp_loaded;
  assign load_pipeline_stages_1_WAYS_TAGS_1_address = ways_1_loadRead_rsp_address;
  assign load_pipeline_stages_1_WAYS_TAGS_1_fault = ways_1_loadRead_rsp_fault;
  assign ways_2_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign ways_2_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[11 : 6];
  assign load_pipeline_stages_1_WAYS_TAGS_2_loaded = ways_2_loadRead_rsp_loaded;
  assign load_pipeline_stages_1_WAYS_TAGS_2_address = ways_2_loadRead_rsp_address;
  assign load_pipeline_stages_1_WAYS_TAGS_2_fault = ways_2_loadRead_rsp_fault;
  assign ways_3_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign ways_3_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[11 : 6];
  assign load_pipeline_stages_1_WAYS_TAGS_3_loaded = ways_3_loadRead_rsp_loaded;
  assign load_pipeline_stages_1_WAYS_TAGS_3_address = ways_3_loadRead_rsp_address;
  assign load_pipeline_stages_1_WAYS_TAGS_3_fault = ways_3_loadRead_rsp_fault;
  assign load_pipeline_stages_2_WAYS_HIT = (|load_pipeline_stages_2_WAYS_HITS);
  assign status_loadRead_cmd_valid = (! (load_pipeline_stages_1_valid && (! load_pipeline_stages_1_ready)));
  assign status_loadRead_cmd_payload = load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[11 : 6];
  assign load_pipeline_stages_1_STATUS_0_dirty = status_loadRead_rsp_0_dirty;
  assign load_pipeline_stages_1_STATUS_1_dirty = status_loadRead_rsp_1_dirty;
  assign load_pipeline_stages_1_STATUS_2_dirty = status_loadRead_rsp_2_dirty;
  assign load_pipeline_stages_1_STATUS_3_dirty = status_loadRead_rsp_3_dirty;
  always @(*) begin
    _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty = load_pipeline_stages_1_STATUS_0_dirty;
    if(when_DataCache_l859) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty = status_writeLast_payload_data_0_dirty;
    end
    if(when_DataCache_l862) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty = status_write_payload_data_0_dirty;
    end
  end

  always @(*) begin
    _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty = load_pipeline_stages_1_STATUS_1_dirty;
    if(when_DataCache_l859) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty = status_writeLast_payload_data_1_dirty;
    end
    if(when_DataCache_l862) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty = status_write_payload_data_1_dirty;
    end
  end

  always @(*) begin
    _zz_load_pipeline_stages_1_STATUS_overloaded_2_dirty = load_pipeline_stages_1_STATUS_2_dirty;
    if(when_DataCache_l859) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_2_dirty = status_writeLast_payload_data_2_dirty;
    end
    if(when_DataCache_l862) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_2_dirty = status_write_payload_data_2_dirty;
    end
  end

  always @(*) begin
    _zz_load_pipeline_stages_1_STATUS_overloaded_3_dirty = load_pipeline_stages_1_STATUS_3_dirty;
    if(when_DataCache_l859) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_3_dirty = status_writeLast_payload_data_3_dirty;
    end
    if(when_DataCache_l862) begin
      _zz_load_pipeline_stages_1_STATUS_overloaded_3_dirty = status_write_payload_data_3_dirty;
    end
  end

  assign when_DataCache_l859 = (status_writeLast_valid && (status_writeLast_payload_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6]));
  assign when_DataCache_l862 = (status_write_valid && (status_write_payload_address == load_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6]));
  assign load_pipeline_stages_1_STATUS_overloaded_0_dirty = _zz_load_pipeline_stages_1_STATUS_overloaded_0_dirty;
  assign load_pipeline_stages_1_STATUS_overloaded_1_dirty = _zz_load_pipeline_stages_1_STATUS_overloaded_1_dirty;
  assign load_pipeline_stages_1_STATUS_overloaded_2_dirty = _zz_load_pipeline_stages_1_STATUS_overloaded_2_dirty;
  assign load_pipeline_stages_1_STATUS_overloaded_3_dirty = _zz_load_pipeline_stages_1_STATUS_overloaded_3_dirty;
  assign load_pipeline_stages_2_REFILL_HITS = {(refill_slots_1_valid && (refill_slots_1_address[31 : 6] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[31 : 6])),(refill_slots_0_valid && (refill_slots_0_address[31 : 6] == load_pipeline_stages_2_ADDRESS_POST_TRANSLATION[31 : 6]))};
  assign load_pipeline_stages_1_LOCKED = (((! load_pipeline_stages_1_UNLOCKED) && io_lock_valid) && (io_lock_address[11 : 6] == load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION[11 : 6]));
  assign load_ctrl_plruLogic_core_evict_logic_0_state = load_ctrl_plruLogic_core_io_context_state_0[0];
  assign load_ctrl_plruLogic_core_evict_sel_0 = (! load_ctrl_plruLogic_core_evict_logic_0_state);
  assign load_ctrl_plruLogic_core_evict_logic_1_stateSel = load_ctrl_plruLogic_core_evict_sel_0;
  assign load_ctrl_plruLogic_core_evict_logic_1_state = load_ctrl_plruLogic_core_io_context_state_1[load_ctrl_plruLogic_core_evict_logic_1_stateSel];
  assign load_ctrl_plruLogic_core_evict_sel_1 = (! load_ctrl_plruLogic_core_evict_logic_1_state);
  assign load_ctrl_plruLogic_core_io_evict_id = {load_ctrl_plruLogic_core_evict_sel_0,load_ctrl_plruLogic_core_evict_sel_1};
  assign load_ctrl_plruLogic_core_io_update_state_0[0] = load_ctrl_plruLogic_core_io_update_id[1];
  assign load_ctrl_plruLogic_core_update_logic_1_sel = load_ctrl_plruLogic_core_io_update_id[1 : 1];
  always @(*) begin
    load_ctrl_plruLogic_core_io_update_state_1 = load_ctrl_plruLogic_core_io_context_state_1;
    load_ctrl_plruLogic_core_io_update_state_1[load_ctrl_plruLogic_core_update_logic_1_sel] = load_ctrl_plruLogic_core_io_update_id[0];
  end

  assign load_ctrl_plruLogic_core_io_context_state_0 = load_pipeline_stages_2_PLRU_0;
  assign load_ctrl_plruLogic_core_io_context_state_1 = load_pipeline_stages_2_PLRU_1;
  always @(*) begin
    load_ctrl_plruLogic_core_io_update_id = 2'bxx;
    if(load_ctrl_startRefill) begin
      load_ctrl_plruLogic_core_io_update_id = load_ctrl_refillWay;
    end
    if(when_DataCache_l1512) begin
      load_ctrl_plruLogic_core_io_update_id = load_ctrl_wayId;
    end
  end

  always @(*) begin
    plru_fromLoad_valid = 1'b0;
    if(load_ctrl_startRefill) begin
      plru_fromLoad_valid = 1'b1;
    end
    if(when_DataCache_l1512) begin
      plru_fromLoad_valid = 1'b1;
    end
  end

  assign plru_fromLoad_payload_address = load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[11 : 6];
  assign plru_fromLoad_payload_data_0 = load_ctrl_plruLogic_core_io_update_state_0;
  assign plru_fromLoad_payload_data_1 = load_ctrl_plruLogic_core_io_update_state_1;
  always @(*) begin
    load_ctrl_reservation_take = 1'b0;
    if(when_DataCache_l1471) begin
      load_ctrl_reservation_take = 1'b1;
    end
  end

  assign load_ctrl_refillWay = load_ctrl_plruLogic_core_io_evict_id;
  assign _zz_refill_push_payload_victim = _zz__zz_refill_push_payload_victim;
  assign load_ctrl_refillWayNeedWriteback = (_zz_load_ctrl_refillWayNeedWriteback && _zz_refill_push_payload_victim);
  assign load_ctrl_refillHit = (|load_pipeline_stages_2_REFILL_HITS);
  assign load_ctrl_refillLoaded = (|({refill_slots_1_loaded,refill_slots_0_loaded} & load_pipeline_stages_2_REFILL_HITS));
  assign load_ctrl_lineBusy = (({(refill_slots_1_valid && (refill_slots_1_address[11 : 6] == load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[11 : 6])),(refill_slots_0_valid && (refill_slots_0_address[11 : 6] == load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION[11 : 6]))} != 2'b00) || 1'b0);
  assign load_ctrl_bankBusy = ((load_pipeline_stages_2_BANK_BUSY_REMAPPED & load_pipeline_stages_2_WAYS_HITS) != 4'b0000);
  assign load_ctrl_waysHitHazard = (|(load_pipeline_stages_2_WAYS_HITS & load_pipeline_stages_2_WAYS_HAZARD_resulting));
  assign load_ctrl_hitUnique = 1'b1;
  assign load_ctrl_uniqueMiss = (load_pipeline_stages_2_NEED_UNIQUE && (! load_ctrl_hitUnique));
  always @(*) begin
    load_pipeline_stages_2_REDO = ((((((! load_pipeline_stages_2_WAYS_HIT) || load_ctrl_waysHitHazard) || load_ctrl_bankBusy) || load_ctrl_refillHit) || load_pipeline_stages_2_LOCKED) || load_ctrl_uniqueMiss);
    if(load_pipeline_stages_2_ABORD) begin
      load_pipeline_stages_2_REDO = 1'b0;
    end
  end

  always @(*) begin
    load_pipeline_stages_2_MISS = ((((! load_pipeline_stages_2_WAYS_HIT) && (! load_ctrl_waysHitHazard)) && (! load_ctrl_refillHit)) && (! load_pipeline_stages_2_LOCKED));
    if(load_pipeline_stages_2_ABORD) begin
      load_pipeline_stages_2_MISS = 1'b0;
    end
  end

  assign load_pipeline_stages_2_FAULT = (|(load_pipeline_stages_2_WAYS_HITS & {load_pipeline_stages_2_WAYS_TAGS_3_fault,{load_pipeline_stages_2_WAYS_TAGS_2_fault,{load_pipeline_stages_2_WAYS_TAGS_1_fault,load_pipeline_stages_2_WAYS_TAGS_0_fault}}}));
  assign load_ctrl_canRefill = (((((! refill_full) && (! load_ctrl_lineBusy)) && load_ctrl_reservation_win) && (! (load_ctrl_refillWayNeedWriteback && writeback_full))) && (! load_pipeline_stages_2_WAYS_HAZARD_resulting[load_ctrl_refillWay]));
  assign load_ctrl_askRefill = ((load_pipeline_stages_2_MISS && load_ctrl_canRefill) && (! load_ctrl_refillHit));
  always @(*) begin
    load_ctrl_askUpgrade = (((! load_pipeline_stages_2_MISS) && load_ctrl_canRefill) && load_ctrl_uniqueMiss);
    if(load_pipeline_stages_2_ABORD) begin
      load_ctrl_askUpgrade = 1'b0;
    end
  end

  assign load_ctrl_startRefill = (load_pipeline_stages_2_valid && load_ctrl_askRefill);
  assign load_ctrl_startUpgrade = (load_pipeline_stages_2_valid && load_ctrl_askUpgrade);
  assign _zz_load_ctrl_wayId = (_zz_load_pipeline_stages_2_CPU_WORD || _zz_load_pipeline_stages_2_CPU_WORD_2);
  assign _zz_load_ctrl_wayId_1 = (_zz_load_pipeline_stages_2_CPU_WORD_1 || _zz_load_pipeline_stages_2_CPU_WORD_2);
  assign load_ctrl_wayId = {_zz_load_ctrl_wayId_1,_zz_load_ctrl_wayId};
  assign when_DataCache_l1471 = (load_ctrl_startRefill || load_ctrl_startUpgrade);
  assign _zz_32 = ({3'd0,1'b1} <<< load_ctrl_refillWay);
  assign when_DataCache_l1512 = ((load_pipeline_stages_2_valid && (! load_pipeline_stages_2_REDO)) && (! load_pipeline_stages_2_MISS));
  assign load_pipeline_stages_2_REFILL_SLOT_FULL = ((load_pipeline_stages_2_MISS && (! load_ctrl_refillHit)) && refill_full);
  assign load_pipeline_stages_2_REFILL_SLOT = (((! load_ctrl_refillLoaded) ? load_pipeline_stages_2_REFILL_HITS : 2'b00) | (load_ctrl_askRefill ? refill_free : 2'b00));
  assign io_load_rsp_valid = load_pipeline_stages_2_valid;
  assign io_load_rsp_payload_data = load_pipeline_stages_2_CPU_WORD;
  assign io_load_rsp_payload_fault = load_pipeline_stages_2_FAULT;
  assign io_load_rsp_payload_redo = load_pipeline_stages_2_REDO;
  assign io_load_rsp_payload_refillSlotAny = load_pipeline_stages_2_REFILL_SLOT_FULL;
  assign io_load_rsp_payload_refillSlot = load_pipeline_stages_2_REFILL_SLOT;
  assign load_pipeline_stages_2_isThrown = load_pipeline_stages_2_throwRequest_DataCache_l1301;
  assign load_pipeline_stages_1_isThrown = load_pipeline_stages_1_throwRequest_DataCache_l1301;
  assign load_pipeline_stages_0_isThrown = load_pipeline_stages_0_throwRequest_DataCache_l1301;
  always @(*) begin
    _zz_load_pipeline_stages_1_valid = load_pipeline_stages_0_valid;
    if(when_Pipeline_l272) begin
      _zz_load_pipeline_stages_1_valid = 1'b0;
    end
  end

  assign load_pipeline_stages_0_ready = 1'b1;
  assign when_Pipeline_l272 = (_zz_load_pipeline_stages_0_throwRequest_DataCache_l1301 != 1'b0);
  always @(*) begin
    _zz_load_pipeline_stages_2_valid = load_pipeline_stages_1_valid;
    if(when_Pipeline_l272_1) begin
      _zz_load_pipeline_stages_2_valid = 1'b0;
    end
  end

  assign load_pipeline_stages_1_ready = 1'b1;
  assign when_Pipeline_l272_1 = (_zz_load_pipeline_stages_1_throwRequest_DataCache_l1301 != 1'b0);
  assign load_pipeline_stages_2_WAYS_HAZARD_resulting = load_pipeline_stages_2_WAYS_HAZARD_overloaded;
  assign store_pipeline_discardAll = 1'b0;
  assign store_pipeline_stages_0_throwRequest_DataCache_l1551 = store_pipeline_discardAll;
  assign store_pipeline_stages_1_throwRequest_DataCache_l1551 = store_pipeline_discardAll;
  assign store_pipeline_stages_2_throwRequest_DataCache_l1551 = store_pipeline_discardAll;
  assign store_pipeline_stages_1_WAYS_HAZARD_overloaded = (store_pipeline_stages_1_WAYS_HAZARD | ((waysWrite_addressLast == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6]) ? waysWrite_maskLast : 4'b0000));
  assign store_pipeline_stages_2_WAYS_HAZARD_overloaded = (store_pipeline_stages_2_WAYS_HAZARD | ((waysWrite_addressLast == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 6]) ? waysWrite_maskLast : 4'b0000));
  assign store_pipeline_stages_0_valid = io_store_cmd_valid;
  assign store_pipeline_stages_0_ADDRESS_POST_TRANSLATION = io_store_cmd_payload_address;
  assign store_pipeline_stages_0_CPU_WORD = io_store_cmd_payload_data;
  assign store_pipeline_stages_0_CPU_MASK = io_store_cmd_payload_mask;
  assign store_pipeline_stages_0_IO = (io_store_cmd_payload_io && (! io_store_cmd_payload_flush));
  assign store_pipeline_stages_0_FLUSH = io_store_cmd_payload_flush;
  assign store_pipeline_stages_0_FLUSH_FREE = io_store_cmd_payload_flushFree;
  assign store_pipeline_stages_0_PREFETCH = io_store_cmd_payload_prefetch;
  assign store_pipeline_stages_0_GENERATION = io_store_cmd_payload_generation;
  assign store_pipeline_stages_0_WAYS_HAZARD = 4'b0000;
  assign io_store_cmd_ready = 1'b1;
  assign _zz_store_pipeline_stages_1_PLRU_0 = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6];
  assign _zz_store_pipeline_stages_1_PLRU_0_1 = _zz_plru_ram_port2;
  assign store_pipeline_stages_1_PLRU_0 = _zz_store_pipeline_stages_1_PLRU_0_1[0 : 0];
  assign store_pipeline_stages_1_PLRU_1 = _zz_store_pipeline_stages_1_PLRU_0_1[2 : 1];
  assign ways_0_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign ways_0_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6];
  assign store_pipeline_stages_1_WAYS_TAGS_0_loaded = ways_0_storeRead_rsp_loaded;
  assign store_pipeline_stages_1_WAYS_TAGS_0_address = ways_0_storeRead_rsp_address;
  assign store_pipeline_stages_1_WAYS_TAGS_0_fault = ways_0_storeRead_rsp_fault;
  always @(*) begin
    store_pipeline_stages_1_WAYS_HITS[0] = (store_pipeline_stages_1_WAYS_TAGS_0_loaded && (store_pipeline_stages_1_WAYS_TAGS_0_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 12]));
    store_pipeline_stages_1_WAYS_HITS[1] = (store_pipeline_stages_1_WAYS_TAGS_1_loaded && (store_pipeline_stages_1_WAYS_TAGS_1_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 12]));
    store_pipeline_stages_1_WAYS_HITS[2] = (store_pipeline_stages_1_WAYS_TAGS_2_loaded && (store_pipeline_stages_1_WAYS_TAGS_2_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 12]));
    store_pipeline_stages_1_WAYS_HITS[3] = (store_pipeline_stages_1_WAYS_TAGS_3_loaded && (store_pipeline_stages_1_WAYS_TAGS_3_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 12]));
  end

  assign ways_1_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign ways_1_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6];
  assign store_pipeline_stages_1_WAYS_TAGS_1_loaded = ways_1_storeRead_rsp_loaded;
  assign store_pipeline_stages_1_WAYS_TAGS_1_address = ways_1_storeRead_rsp_address;
  assign store_pipeline_stages_1_WAYS_TAGS_1_fault = ways_1_storeRead_rsp_fault;
  assign ways_2_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign ways_2_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6];
  assign store_pipeline_stages_1_WAYS_TAGS_2_loaded = ways_2_storeRead_rsp_loaded;
  assign store_pipeline_stages_1_WAYS_TAGS_2_address = ways_2_storeRead_rsp_address;
  assign store_pipeline_stages_1_WAYS_TAGS_2_fault = ways_2_storeRead_rsp_fault;
  assign ways_3_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign ways_3_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6];
  assign store_pipeline_stages_1_WAYS_TAGS_3_loaded = ways_3_storeRead_rsp_loaded;
  assign store_pipeline_stages_1_WAYS_TAGS_3_address = ways_3_storeRead_rsp_address;
  assign store_pipeline_stages_1_WAYS_TAGS_3_fault = ways_3_storeRead_rsp_fault;
  assign store_pipeline_stages_1_WAYS_HIT = (|store_pipeline_stages_1_WAYS_HITS);
  assign status_storeRead_cmd_valid = (! (store_pipeline_stages_1_valid && (! store_pipeline_stages_1_ready)));
  assign status_storeRead_cmd_payload = store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6];
  assign store_pipeline_stages_1_STATUS_0_dirty = status_storeRead_rsp_0_dirty;
  assign store_pipeline_stages_1_STATUS_1_dirty = status_storeRead_rsp_1_dirty;
  assign store_pipeline_stages_1_STATUS_2_dirty = status_storeRead_rsp_2_dirty;
  assign store_pipeline_stages_1_STATUS_3_dirty = status_storeRead_rsp_3_dirty;
  always @(*) begin
    _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty = store_pipeline_stages_1_STATUS_0_dirty;
    if(when_DataCache_l859_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty = status_writeLast_payload_data_0_dirty;
    end
    if(when_DataCache_l862_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty = status_write_payload_data_0_dirty;
    end
  end

  always @(*) begin
    _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty = store_pipeline_stages_1_STATUS_1_dirty;
    if(when_DataCache_l859_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty = status_writeLast_payload_data_1_dirty;
    end
    if(when_DataCache_l862_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty = status_write_payload_data_1_dirty;
    end
  end

  always @(*) begin
    _zz_store_pipeline_stages_1_STATUS_overloaded_2_dirty = store_pipeline_stages_1_STATUS_2_dirty;
    if(when_DataCache_l859_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_2_dirty = status_writeLast_payload_data_2_dirty;
    end
    if(when_DataCache_l862_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_2_dirty = status_write_payload_data_2_dirty;
    end
  end

  always @(*) begin
    _zz_store_pipeline_stages_1_STATUS_overloaded_3_dirty = store_pipeline_stages_1_STATUS_3_dirty;
    if(when_DataCache_l859_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_3_dirty = status_writeLast_payload_data_3_dirty;
    end
    if(when_DataCache_l862_1) begin
      _zz_store_pipeline_stages_1_STATUS_overloaded_3_dirty = status_write_payload_data_3_dirty;
    end
  end

  assign when_DataCache_l859_1 = (status_writeLast_valid && (status_writeLast_payload_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6]));
  assign when_DataCache_l862_1 = (status_write_valid && (status_write_payload_address == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[11 : 6]));
  assign store_pipeline_stages_1_STATUS_overloaded_0_dirty = _zz_store_pipeline_stages_1_STATUS_overloaded_0_dirty;
  assign store_pipeline_stages_1_STATUS_overloaded_1_dirty = _zz_store_pipeline_stages_1_STATUS_overloaded_1_dirty;
  assign store_pipeline_stages_1_STATUS_overloaded_2_dirty = _zz_store_pipeline_stages_1_STATUS_overloaded_2_dirty;
  assign store_pipeline_stages_1_STATUS_overloaded_3_dirty = _zz_store_pipeline_stages_1_STATUS_overloaded_3_dirty;
  always @(*) begin
    store_pipeline_stages_1_REFILL_HITS_EARLY = {(refill_slots_1_valid && (refill_slots_1_address[31 : 6] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 6])),(refill_slots_0_valid && (refill_slots_0_address[31 : 6] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 6]))};
    if(store_refillCheckEarly_refillPushHit) begin
      if(_zz_27) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[0] = 1'b1;
      end
      if(_zz_28) begin
        store_pipeline_stages_1_REFILL_HITS_EARLY[1] = 1'b1;
      end
    end
  end

  assign store_refillCheckEarly_refillPushHit = (refill_push_valid && (refill_push_payload_address[31 : 6] == store_pipeline_stages_1_ADDRESS_POST_TRANSLATION[31 : 6]));
  assign store_pipeline_stages_2_REFILL_HITS = (store_pipeline_stages_2_REFILL_HITS_EARLY & {refill_slots_1_valid,refill_slots_0_valid});
  assign store_pipeline_stages_2_PROBE = 1'b0;
  assign store_ctrl_plruLogic_core_evict_logic_0_state = store_ctrl_plruLogic_core_io_context_state_0[0];
  assign store_ctrl_plruLogic_core_evict_sel_0 = (! store_ctrl_plruLogic_core_evict_logic_0_state);
  assign store_ctrl_plruLogic_core_evict_logic_1_stateSel = store_ctrl_plruLogic_core_evict_sel_0;
  assign store_ctrl_plruLogic_core_evict_logic_1_state = store_ctrl_plruLogic_core_io_context_state_1[store_ctrl_plruLogic_core_evict_logic_1_stateSel];
  assign store_ctrl_plruLogic_core_evict_sel_1 = (! store_ctrl_plruLogic_core_evict_logic_1_state);
  assign store_ctrl_plruLogic_core_io_evict_id = {store_ctrl_plruLogic_core_evict_sel_0,store_ctrl_plruLogic_core_evict_sel_1};
  assign store_ctrl_plruLogic_core_io_update_state_0[0] = store_ctrl_plruLogic_core_io_update_id[1];
  assign store_ctrl_plruLogic_core_update_logic_1_sel = store_ctrl_plruLogic_core_io_update_id[1 : 1];
  always @(*) begin
    store_ctrl_plruLogic_core_io_update_state_1 = store_ctrl_plruLogic_core_io_context_state_1;
    store_ctrl_plruLogic_core_io_update_state_1[store_ctrl_plruLogic_core_update_logic_1_sel] = store_ctrl_plruLogic_core_io_update_id[0];
  end

  assign store_ctrl_plruLogic_core_io_context_state_0 = store_pipeline_stages_2_PLRU_0;
  assign store_ctrl_plruLogic_core_io_context_state_1 = store_pipeline_stages_2_PLRU_1;
  always @(*) begin
    store_ctrl_plruLogic_core_io_update_id = 2'bxx;
    if(store_ctrl_startRefill) begin
      store_ctrl_plruLogic_core_io_update_id = store_ctrl_refillWay;
    end
    if(store_ctrl_writeCache) begin
      store_ctrl_plruLogic_core_io_update_id = store_ctrl_wayId;
    end
  end

  always @(*) begin
    plru_fromStore_valid = 1'b0;
    if(store_ctrl_startRefill) begin
      plru_fromStore_valid = 1'b1;
    end
    if(store_ctrl_writeCache) begin
      plru_fromStore_valid = 1'b1;
    end
  end

  assign plru_fromStore_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 6];
  assign plru_fromStore_payload_data_0 = store_ctrl_plruLogic_core_io_update_state_0;
  assign plru_fromStore_payload_data_1 = store_ctrl_plruLogic_core_io_update_state_1;
  assign store_pipeline_stages_2_GENERATION_OK = (((store_pipeline_stages_2_GENERATION == store_target) || store_pipeline_stages_2_PREFETCH) || store_pipeline_stages_2_PROBE);
  always @(*) begin
    store_ctrl_reservation_take = 1'b0;
    if(when_DataCache_l1725) begin
      store_ctrl_reservation_take = 1'b1;
    end
  end

  assign store_ctrl_replacedWay = store_ctrl_plruLogic_core_io_evict_id;
  assign store_ctrl_replacedWayNeedWriteback = (_zz_store_ctrl_replacedWayNeedWriteback && _zz_store_ctrl_replacedWayNeedWriteback_1);
  assign store_ctrl_refillHit = (|(store_pipeline_stages_2_REFILL_HITS & {refill_slots_1_valid,refill_slots_0_valid}));
  assign store_ctrl_lineBusy = (({(refill_slots_1_valid && (refill_slots_1_address[11 : 6] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 6])),(refill_slots_0_valid && (refill_slots_0_address[11 : 6] == store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[11 : 6]))} != 2'b00) || 1'b0);
  assign store_ctrl_waysHitHazard = (|(store_pipeline_stages_2_WAYS_HITS & store_pipeline_stages_2_WAYS_HAZARD_resulting));
  assign store_ctrl_wasClean = (! (|({store_pipeline_stages_2_STATUS_3_dirty,{store_pipeline_stages_2_STATUS_2_dirty,{store_pipeline_stages_2_STATUS_1_dirty,store_pipeline_stages_2_STATUS_0_dirty}}} & store_pipeline_stages_2_WAYS_HITS)));
  assign store_ctrl_bankBusy = ((((! store_pipeline_stages_2_FLUSH) && (! store_pipeline_stages_2_PREFETCH)) && (! store_pipeline_stages_2_PROBE)) && (|(store_pipeline_stages_2_WAYS_HITS & refill_read_bankWriteNotif)));
  assign store_ctrl_hitUnique = 1'b1;
  assign store_ctrl_hitFault = (|(store_pipeline_stages_2_WAYS_HITS & {store_pipeline_stages_2_WAYS_TAGS_3_fault,{store_pipeline_stages_2_WAYS_TAGS_2_fault,{store_pipeline_stages_2_WAYS_TAGS_1_fault,store_pipeline_stages_2_WAYS_TAGS_0_fault}}}));
  always @(*) begin
    store_ctrl_refillWay = store_ctrl_replacedWay;
    if(when_DataCache_l1705) begin
      store_ctrl_refillWay = store_ctrl_wayId;
    end
  end

  always @(*) begin
    store_pipeline_stages_2_REDO = (((((store_pipeline_stages_2_MISS || store_ctrl_waysHitHazard) || store_ctrl_bankBusy) || store_ctrl_refillHit) || (store_ctrl_wasClean && (! store_ctrl_reservation_win))) || (! store_ctrl_hitUnique));
    if(store_pipeline_stages_2_FLUSH) begin
      store_pipeline_stages_2_REDO = (store_ctrl_needFlush || (|store_pipeline_stages_2_WAYS_HAZARD_resulting));
    end
    if(store_pipeline_stages_2_IO) begin
      store_pipeline_stages_2_REDO = 1'b0;
    end
  end

  always @(*) begin
    store_pipeline_stages_2_MISS = (((! store_pipeline_stages_2_WAYS_HIT) && (! store_ctrl_waysHitHazard)) && (! store_ctrl_refillHit));
    if(store_pipeline_stages_2_IO) begin
      store_pipeline_stages_2_MISS = 1'b0;
    end
  end

  assign store_ctrl_canRefill = (((((! refill_full) && (! store_ctrl_lineBusy)) && (! load_ctrl_startRefill)) && store_ctrl_reservation_win) && (! store_pipeline_stages_2_WAYS_HAZARD_resulting[store_ctrl_refillWay]));
  assign store_ctrl_askRefill = (((store_pipeline_stages_2_MISS && store_ctrl_canRefill) && (! store_ctrl_refillHit)) && (! (store_ctrl_replacedWayNeedWriteback && writeback_full)));
  assign store_ctrl_askUpgrade = (((! store_pipeline_stages_2_MISS) && store_ctrl_canRefill) && (! store_ctrl_hitUnique));
  always @(*) begin
    store_ctrl_startRefill = ((store_pipeline_stages_2_valid && store_pipeline_stages_2_GENERATION_OK) && store_ctrl_askRefill);
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_startRefill = 1'b0;
    end
  end

  always @(*) begin
    store_ctrl_startUpgrade = ((store_pipeline_stages_2_valid && store_pipeline_stages_2_GENERATION_OK) && store_ctrl_askUpgrade);
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_startUpgrade = 1'b0;
    end
    if(store_pipeline_stages_2_IO) begin
      store_ctrl_startUpgrade = 1'b0;
    end
  end

  assign store_pipeline_stages_2_REFILL_SLOT_FULL = ((store_pipeline_stages_2_MISS && (! store_ctrl_refillHit)) && refill_full);
  assign store_pipeline_stages_2_REFILL_SLOT = ((store_ctrl_askRefill || store_ctrl_askUpgrade) ? refill_free : 2'b00);
  always @(*) begin
    store_ctrl_writeCache = ((((store_pipeline_stages_2_valid && store_pipeline_stages_2_GENERATION_OK) && (! store_pipeline_stages_2_REDO)) && (! store_pipeline_stages_2_PREFETCH)) && (! store_pipeline_stages_2_PROBE));
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_writeCache = 1'b0;
    end
    if(store_pipeline_stages_2_IO) begin
      store_ctrl_writeCache = 1'b0;
    end
  end

  always @(*) begin
    store_ctrl_setDirty = (store_ctrl_writeCache && store_ctrl_wasClean);
    if(store_pipeline_stages_2_FLUSH) begin
      store_ctrl_setDirty = 1'b0;
    end
    if(store_pipeline_stages_2_IO) begin
      store_ctrl_setDirty = 1'b0;
    end
  end

  assign _zz_store_ctrl_wayId = store_pipeline_stages_2_WAYS_HITS[1];
  assign _zz_store_ctrl_wayId_1 = store_pipeline_stages_2_WAYS_HITS[2];
  assign _zz_store_ctrl_wayId_2 = store_pipeline_stages_2_WAYS_HITS[3];
  assign _zz_store_ctrl_wayId_3 = (_zz_store_ctrl_wayId || _zz_store_ctrl_wayId_2);
  assign _zz_store_ctrl_wayId_4 = (_zz_store_ctrl_wayId_1 || _zz_store_ctrl_wayId_2);
  assign store_ctrl_wayId = {_zz_store_ctrl_wayId_4,_zz_store_ctrl_wayId_3};
  assign store_ctrl_needFlushs = ({store_pipeline_stages_2_WAYS_TAGS_3_loaded,{store_pipeline_stages_2_WAYS_TAGS_2_loaded,{store_pipeline_stages_2_WAYS_TAGS_1_loaded,store_pipeline_stages_2_WAYS_TAGS_0_loaded}}} & {store_pipeline_stages_2_STATUS_3_dirty,{store_pipeline_stages_2_STATUS_2_dirty,{store_pipeline_stages_2_STATUS_1_dirty,store_pipeline_stages_2_STATUS_0_dirty}}});
  assign _zz_store_ctrl_needFlushs_bools_0 = store_ctrl_needFlushs;
  assign store_ctrl_needFlushs_bools_0 = _zz_store_ctrl_needFlushs_bools_0[0];
  assign store_ctrl_needFlushs_bools_1 = _zz_store_ctrl_needFlushs_bools_0[1];
  assign store_ctrl_needFlushs_bools_2 = _zz_store_ctrl_needFlushs_bools_0[2];
  assign store_ctrl_needFlushs_bools_3 = _zz_store_ctrl_needFlushs_bools_0[3];
  always @(*) begin
    _zz_store_ctrl_needFlushOh[0] = (store_ctrl_needFlushs_bools_0 && (! 1'b0));
    _zz_store_ctrl_needFlushOh[1] = (store_ctrl_needFlushs_bools_1 && (! store_ctrl_needFlushs_bools_0));
    _zz_store_ctrl_needFlushOh[2] = (store_ctrl_needFlushs_bools_2 && (! store_ctrl_needFlushs_range_0_to_1));
    _zz_store_ctrl_needFlushOh[3] = (store_ctrl_needFlushs_bools_3 && (! store_ctrl_needFlushs_range_0_to_2));
  end

  assign store_ctrl_needFlushs_range_0_to_1 = ({store_ctrl_needFlushs_bools_1,store_ctrl_needFlushs_bools_0} != 2'b00);
  assign store_ctrl_needFlushs_range_0_to_2 = ({store_ctrl_needFlushs_bools_2,{store_ctrl_needFlushs_bools_1,store_ctrl_needFlushs_bools_0}} != 3'b000);
  assign store_ctrl_needFlushOh = _zz_store_ctrl_needFlushOh;
  assign _zz_34 = store_ctrl_needFlushOh[0];
  assign _zz_store_ctrl_needFlushSel = store_ctrl_needFlushOh[1];
  assign _zz_store_ctrl_needFlushSel_1 = store_ctrl_needFlushOh[2];
  assign _zz_store_ctrl_needFlushSel_2 = store_ctrl_needFlushOh[3];
  assign _zz_store_ctrl_needFlushSel_3 = (_zz_store_ctrl_needFlushSel || _zz_store_ctrl_needFlushSel_2);
  assign _zz_store_ctrl_needFlushSel_4 = (_zz_store_ctrl_needFlushSel_1 || _zz_store_ctrl_needFlushSel_2);
  assign store_ctrl_needFlushSel = {_zz_store_ctrl_needFlushSel_4,_zz_store_ctrl_needFlushSel_3};
  assign store_ctrl_needFlush = (|store_ctrl_needFlushs);
  assign store_ctrl_canFlush = (((store_ctrl_reservation_win && (! writeback_full)) && (! ({refill_slots_1_valid,refill_slots_0_valid} != 2'b00))) && (! (|store_pipeline_stages_2_WAYS_HAZARD_resulting)));
  assign store_ctrl_startFlush = ((((store_pipeline_stages_2_valid && store_pipeline_stages_2_FLUSH) && store_pipeline_stages_2_GENERATION_OK) && store_ctrl_needFlush) && store_ctrl_canFlush);
  assign when_DataCache_l1705 = ((! store_pipeline_stages_2_MISS) && (! store_ctrl_hitUnique));
  assign when_DataCache_l1725 = (((store_ctrl_startRefill || store_ctrl_startUpgrade) || store_ctrl_setDirty) || store_ctrl_startFlush);
  assign when_DataCache_l1732 = (store_ctrl_startRefill || store_ctrl_startFlush);
  assign when_DataCache_l1750 = (store_ctrl_startRefill || store_ctrl_startUpgrade);
  assign when_DataCache_l1774 = store_pipeline_stages_2_WAYS_HITS[0];
  assign _zz_35 = ({1'd0,1'b1} <<< store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[2 : 2]);
  assign when_DataCache_l1774_1 = store_pipeline_stages_2_WAYS_HITS[1];
  assign _zz_36 = ({1'd0,1'b1} <<< store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[2 : 2]);
  assign when_DataCache_l1774_2 = store_pipeline_stages_2_WAYS_HITS[2];
  assign _zz_37 = ({1'd0,1'b1} <<< store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[2 : 2]);
  assign when_DataCache_l1774_3 = store_pipeline_stages_2_WAYS_HITS[3];
  assign _zz_38 = ({1'd0,1'b1} <<< store_pipeline_stages_2_ADDRESS_POST_TRANSLATION[2 : 2]);
  assign when_DataCache_l1804 = ((((store_pipeline_stages_2_valid && store_pipeline_stages_2_REDO) && store_pipeline_stages_2_GENERATION_OK) && (! store_pipeline_stages_2_PREFETCH)) && (! store_pipeline_stages_2_PROBE));
  assign io_store_rsp_valid = (store_pipeline_stages_2_valid && (! store_pipeline_stages_2_PROBE));
  assign io_store_rsp_payload_generationKo = (! store_pipeline_stages_2_GENERATION_OK);
  assign io_store_rsp_payload_fault = 1'b0;
  assign io_store_rsp_payload_redo = store_pipeline_stages_2_REDO;
  assign io_store_rsp_payload_refillSlotAny = store_pipeline_stages_2_REFILL_SLOT_FULL;
  assign io_store_rsp_payload_refillSlot = store_pipeline_stages_2_REFILL_SLOT;
  assign io_store_rsp_payload_flush = store_pipeline_stages_2_FLUSH;
  assign io_store_rsp_payload_prefetch = store_pipeline_stages_2_PREFETCH;
  assign io_store_rsp_payload_address = store_pipeline_stages_2_ADDRESS_POST_TRANSLATION;
  assign io_store_rsp_payload_io = store_pipeline_stages_2_IO;
  assign store_pipeline_stages_2_isThrown = store_pipeline_stages_2_throwRequest_DataCache_l1551;
  assign store_pipeline_stages_1_isThrown = store_pipeline_stages_1_throwRequest_DataCache_l1551;
  assign store_pipeline_stages_0_isThrown = store_pipeline_stages_0_throwRequest_DataCache_l1551;
  always @(*) begin
    _zz_store_pipeline_stages_1_valid = store_pipeline_stages_0_valid;
    if(when_Pipeline_l272_2) begin
      _zz_store_pipeline_stages_1_valid = 1'b0;
    end
  end

  assign when_Pipeline_l272_2 = (store_pipeline_discardAll != 1'b0);
  always @(*) begin
    _zz_store_pipeline_stages_2_valid = store_pipeline_stages_1_valid;
    if(when_Pipeline_l272_3) begin
      _zz_store_pipeline_stages_2_valid = 1'b0;
    end
  end

  assign store_pipeline_stages_1_ready = 1'b1;
  assign when_Pipeline_l272_3 = (store_pipeline_discardAll != 1'b0);
  assign store_pipeline_stages_2_WAYS_HAZARD_resulting = store_pipeline_stages_2_WAYS_HAZARD_overloaded;
  assign io_refillEvent = refill_push_valid;
  assign io_writebackEvent = writeback_push_valid;
  assign io_tagEvent = (|waysWrite_mask);
  assign invalidate_reservation_win = (! 1'b0);
  assign refill_read_reservation_win = (! 1'b0);
  assign load_ctrl_reservation_win = (! ({refill_read_reservation_take,invalidate_reservation_take} != 2'b00));
  assign store_ctrl_reservation_win = (! ({load_ctrl_reservation_take,{refill_read_reservation_take,invalidate_reservation_take}} != 3'b000));
  always @(*) begin
    _zz_banks_0_read_rsp = _zz_banks_0_mem_port1;
    if(when_MultiportRam_l328) begin
      if(_zz_39[0]) begin
        _zz_banks_0_read_rsp[7 : 0] = 8'bxxxxxxxx;
      end
      if(_zz_39[1]) begin
        _zz_banks_0_read_rsp[15 : 8] = 8'bxxxxxxxx;
      end
      if(_zz_39[2]) begin
        _zz_banks_0_read_rsp[23 : 16] = 8'bxxxxxxxx;
      end
      if(_zz_39[3]) begin
        _zz_banks_0_read_rsp[31 : 24] = 8'bxxxxxxxx;
      end
      if(_zz_39[4]) begin
        _zz_banks_0_read_rsp[39 : 32] = 8'bxxxxxxxx;
      end
      if(_zz_39[5]) begin
        _zz_banks_0_read_rsp[47 : 40] = 8'bxxxxxxxx;
      end
      if(_zz_39[6]) begin
        _zz_banks_0_read_rsp[55 : 48] = 8'bxxxxxxxx;
      end
      if(_zz_39[7]) begin
        _zz_banks_0_read_rsp[63 : 56] = 8'bxxxxxxxx;
      end
    end
  end

  always @(*) begin
    _zz_banks_1_read_rsp = _zz_banks_1_mem_port1;
    if(when_MultiportRam_l328_1) begin
      if(_zz_40[0]) begin
        _zz_banks_1_read_rsp[7 : 0] = 8'bxxxxxxxx;
      end
      if(_zz_40[1]) begin
        _zz_banks_1_read_rsp[15 : 8] = 8'bxxxxxxxx;
      end
      if(_zz_40[2]) begin
        _zz_banks_1_read_rsp[23 : 16] = 8'bxxxxxxxx;
      end
      if(_zz_40[3]) begin
        _zz_banks_1_read_rsp[31 : 24] = 8'bxxxxxxxx;
      end
      if(_zz_40[4]) begin
        _zz_banks_1_read_rsp[39 : 32] = 8'bxxxxxxxx;
      end
      if(_zz_40[5]) begin
        _zz_banks_1_read_rsp[47 : 40] = 8'bxxxxxxxx;
      end
      if(_zz_40[6]) begin
        _zz_banks_1_read_rsp[55 : 48] = 8'bxxxxxxxx;
      end
      if(_zz_40[7]) begin
        _zz_banks_1_read_rsp[63 : 56] = 8'bxxxxxxxx;
      end
    end
  end

  always @(*) begin
    _zz_banks_2_read_rsp = _zz_banks_2_mem_port1;
    if(when_MultiportRam_l328_2) begin
      if(_zz_41[0]) begin
        _zz_banks_2_read_rsp[7 : 0] = 8'bxxxxxxxx;
      end
      if(_zz_41[1]) begin
        _zz_banks_2_read_rsp[15 : 8] = 8'bxxxxxxxx;
      end
      if(_zz_41[2]) begin
        _zz_banks_2_read_rsp[23 : 16] = 8'bxxxxxxxx;
      end
      if(_zz_41[3]) begin
        _zz_banks_2_read_rsp[31 : 24] = 8'bxxxxxxxx;
      end
      if(_zz_41[4]) begin
        _zz_banks_2_read_rsp[39 : 32] = 8'bxxxxxxxx;
      end
      if(_zz_41[5]) begin
        _zz_banks_2_read_rsp[47 : 40] = 8'bxxxxxxxx;
      end
      if(_zz_41[6]) begin
        _zz_banks_2_read_rsp[55 : 48] = 8'bxxxxxxxx;
      end
      if(_zz_41[7]) begin
        _zz_banks_2_read_rsp[63 : 56] = 8'bxxxxxxxx;
      end
    end
  end

  always @(*) begin
    _zz_banks_3_read_rsp = _zz_banks_3_mem_port1;
    if(when_MultiportRam_l328_3) begin
      if(_zz_42[0]) begin
        _zz_banks_3_read_rsp[7 : 0] = 8'bxxxxxxxx;
      end
      if(_zz_42[1]) begin
        _zz_banks_3_read_rsp[15 : 8] = 8'bxxxxxxxx;
      end
      if(_zz_42[2]) begin
        _zz_banks_3_read_rsp[23 : 16] = 8'bxxxxxxxx;
      end
      if(_zz_42[3]) begin
        _zz_banks_3_read_rsp[31 : 24] = 8'bxxxxxxxx;
      end
      if(_zz_42[4]) begin
        _zz_banks_3_read_rsp[39 : 32] = 8'bxxxxxxxx;
      end
      if(_zz_42[5]) begin
        _zz_banks_3_read_rsp[47 : 40] = 8'bxxxxxxxx;
      end
      if(_zz_42[6]) begin
        _zz_banks_3_read_rsp[55 : 48] = 8'bxxxxxxxx;
      end
      if(_zz_42[7]) begin
        _zz_banks_3_read_rsp[63 : 56] = 8'bxxxxxxxx;
      end
    end
  end

  always @(*) begin
    _zz_writeback_write_word = _zz_writeback_victimBuffer_port1;
    if(when_MultiportRam_l328_4) begin
      _zz_writeback_write_word = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    end
  end

  always @(posedge clk) begin
    waysWrite_maskLast <= waysWrite_mask;
    waysWrite_addressLast <= waysWrite_address;
    status_writeLast_payload_address <= status_write_payload_address;
    status_writeLast_payload_data_0_dirty <= status_write_payload_data_0_dirty;
    status_writeLast_payload_data_1_dirty <= status_write_payload_data_1_dirty;
    status_writeLast_payload_data_2_dirty <= status_write_payload_data_2_dirty;
    status_writeLast_payload_data_3_dirty <= status_write_payload_data_3_dirty;
    refill_slots_0_loadedCounter <= (refill_slots_0_loadedCounter + (refill_slots_0_loaded && (! refill_slots_0_loadedDone)));
    refill_slots_1_loadedCounter <= (refill_slots_1_loadedCounter + (refill_slots_1_loaded && (! refill_slots_1_loadedDone)));
    if(refill_push_valid) begin
      if(when_DataCache_l960) begin
        refill_slots_0_address <= refill_push_payload_address;
        refill_slots_0_way <= refill_push_payload_way;
        refill_slots_0_cmdSent <= 1'b0;
        refill_slots_0_priority <= 1'b1;
        refill_slots_0_loaded <= 1'b0;
        refill_slots_0_loadedCounter <= 1'b0;
        refill_slots_0_victim <= refill_push_payload_victim;
        refill_slots_0_writebackHazards <= 2'b00;
      end else begin
        if(_zz_28) begin
          refill_slots_0_priority[0] <= 1'b0;
        end
      end
    end
    if(refill_push_valid) begin
      if(when_DataCache_l960_1) begin
        refill_slots_1_address <= refill_push_payload_address;
        refill_slots_1_way <= refill_push_payload_way;
        refill_slots_1_cmdSent <= 1'b0;
        refill_slots_1_priority <= 1'b1;
        refill_slots_1_loaded <= 1'b0;
        refill_slots_1_loadedCounter <= 1'b0;
        refill_slots_1_victim <= refill_push_payload_victim;
        refill_slots_1_writebackHazards <= 2'b00;
      end else begin
        if(_zz_27) begin
          refill_slots_1_priority[0] <= 1'b0;
        end
      end
    end
    if(refill_read_arbiter_oh[0]) begin
      refill_slots_0_writebackHazards <= refill_read_writebackHazards;
      if(when_DataCache_l997) begin
        refill_slots_0_cmdSent <= 1'b1;
      end
    end
    if(_zz_refill_read_arbiter_sel) begin
      refill_slots_1_writebackHazards <= refill_read_writebackHazards;
      if(when_DataCache_l997_1) begin
        refill_slots_1_cmdSent <= 1'b1;
      end
    end
    if(io_mem_read_rsp_valid) begin
      if(when_DataCache_l1036) begin
        case(io_mem_read_rsp_payload_id)
          1'b0 : begin
            refill_slots_0_loaded <= 1'b1;
          end
          default : begin
            refill_slots_1_loaded <= 1'b1;
          end
        endcase
      end
    end
    if(writeback_slots_0_fire) begin
      refill_slots_0_writebackHazards[0] <= 1'b0;
      refill_slots_1_writebackHazards[0] <= 1'b0;
    end
    if(writeback_slots_1_fire) begin
      refill_slots_0_writebackHazards[1] <= 1'b0;
      refill_slots_1_writebackHazards[1] <= 1'b0;
    end
    if(writeback_push_valid) begin
      if(when_DataCache_l1127) begin
        writeback_slots_0_address <= writeback_push_payload_address;
        writeback_slots_0_way <= writeback_push_payload_way;
        writeback_slots_0_writeCmdDone <= 1'b0;
        writeback_slots_0_priority <= 1'b1;
        writeback_slots_0_readCmdDone <= 1'b0;
        writeback_slots_0_readRspDone <= 1'b0;
        writeback_slots_0_victimBufferReady <= 1'b0;
      end else begin
        if(writeback_free[1]) begin
          writeback_slots_0_priority[0] <= 1'b0;
        end
      end
    end
    if(writeback_push_valid) begin
      if(when_DataCache_l1127_1) begin
        writeback_slots_1_address <= writeback_push_payload_address;
        writeback_slots_1_way <= writeback_push_payload_way;
        writeback_slots_1_writeCmdDone <= 1'b0;
        writeback_slots_1_priority <= 1'b1;
        writeback_slots_1_readCmdDone <= 1'b0;
        writeback_slots_1_readRspDone <= 1'b0;
        writeback_slots_1_victimBufferReady <= 1'b0;
      end else begin
        if(writeback_free[0]) begin
          writeback_slots_1_priority[0] <= 1'b0;
        end
      end
    end
    if(when_DataCache_l1174) begin
      if(writeback_read_arbiter_oh[0]) begin
        writeback_slots_0_readCmdDone <= 1'b1;
      end
      if(_zz_writeback_read_arbiter_sel) begin
        writeback_slots_1_readCmdDone <= 1'b1;
      end
    end
    if(writeback_read_slotRead_valid) begin
      refill_slots_0_victim[writeback_read_slotRead_payload_id] <= 1'b0;
      refill_slots_1_victim[writeback_read_slotRead_payload_id] <= 1'b0;
    end
    writeback_read_slotReadLast_payload_id <= writeback_read_slotRead_payload_id;
    writeback_read_slotReadLast_payload_last <= writeback_read_slotRead_payload_last;
    writeback_read_slotReadLast_payload_wordIndex <= writeback_read_slotRead_payload_wordIndex;
    writeback_read_slotReadLast_payload_way <= writeback_read_slotRead_payload_way;
    if(writeback_read_slotReadLast_valid) begin
      case(writeback_read_slotReadLast_payload_id)
        1'b0 : begin
          writeback_slots_0_victimBufferReady <= 1'b1;
        end
        default : begin
          writeback_slots_1_victimBufferReady <= 1'b1;
        end
      endcase
      if(writeback_read_slotReadLast_payload_last) begin
        case(writeback_read_slotReadLast_payload_id)
          1'b0 : begin
            writeback_slots_0_readRspDone <= 1'b1;
          end
          default : begin
            writeback_slots_1_readRspDone <= 1'b1;
          end
        endcase
      end
    end
    if(when_DataCache_l1252) begin
      if(writeback_write_arbiter_oh[0]) begin
        writeback_slots_0_writeCmdDone <= 1'b1;
      end
      if(_zz_writeback_write_arbiter_sel) begin
        writeback_slots_1_writeCmdDone <= 1'b1;
      end
    end
    if(writeback_write_bufferRead_ready) begin
      writeback_write_bufferRead_rData_id <= writeback_write_bufferRead_payload_id;
      writeback_write_bufferRead_rData_address <= writeback_write_bufferRead_payload_address;
      writeback_write_bufferRead_rData_last <= writeback_write_bufferRead_payload_last;
    end
    load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION <= load_pipeline_stages_0_ADDRESS_PRE_TRANSLATION;
    load_pipeline_stages_1_WAYS_HAZARD <= load_pipeline_stages_0_WAYS_HAZARD;
    load_pipeline_stages_1_UNLOCKED <= load_pipeline_stages_0_UNLOCKED;
    load_pipeline_stages_1_NEED_UNIQUE <= load_pipeline_stages_0_NEED_UNIQUE;
    load_pipeline_stages_1_BANK_BUSY <= load_pipeline_stages_0_BANK_BUSY_overloaded;
    load_pipeline_stages_2_WAYS_HAZARD <= load_pipeline_stages_1_WAYS_HAZARD_overloaded;
    load_pipeline_stages_2_ADDRESS_PRE_TRANSLATION <= load_pipeline_stages_1_ADDRESS_PRE_TRANSLATION;
    load_pipeline_stages_2_BANK_BUSY_REMAPPED <= load_pipeline_stages_1_BANK_BUSY_REMAPPED;
    load_pipeline_stages_2_BANKS_MUXES_0 <= load_pipeline_stages_1_BANKS_MUXES_0;
    load_pipeline_stages_2_BANKS_MUXES_1 <= load_pipeline_stages_1_BANKS_MUXES_1;
    load_pipeline_stages_2_BANKS_MUXES_2 <= load_pipeline_stages_1_BANKS_MUXES_2;
    load_pipeline_stages_2_BANKS_MUXES_3 <= load_pipeline_stages_1_BANKS_MUXES_3;
    load_pipeline_stages_2_ADDRESS_POST_TRANSLATION <= load_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
    load_pipeline_stages_2_ABORD <= load_pipeline_stages_1_ABORD;
    load_pipeline_stages_2_PLRU_0 <= load_pipeline_stages_1_PLRU_0;
    load_pipeline_stages_2_PLRU_1 <= load_pipeline_stages_1_PLRU_1;
    load_pipeline_stages_2_WAYS_TAGS_0_loaded <= load_pipeline_stages_1_WAYS_TAGS_0_loaded;
    load_pipeline_stages_2_WAYS_TAGS_0_address <= load_pipeline_stages_1_WAYS_TAGS_0_address;
    load_pipeline_stages_2_WAYS_TAGS_0_fault <= load_pipeline_stages_1_WAYS_TAGS_0_fault;
    load_pipeline_stages_2_WAYS_TAGS_1_loaded <= load_pipeline_stages_1_WAYS_TAGS_1_loaded;
    load_pipeline_stages_2_WAYS_TAGS_1_address <= load_pipeline_stages_1_WAYS_TAGS_1_address;
    load_pipeline_stages_2_WAYS_TAGS_1_fault <= load_pipeline_stages_1_WAYS_TAGS_1_fault;
    load_pipeline_stages_2_WAYS_TAGS_2_loaded <= load_pipeline_stages_1_WAYS_TAGS_2_loaded;
    load_pipeline_stages_2_WAYS_TAGS_2_address <= load_pipeline_stages_1_WAYS_TAGS_2_address;
    load_pipeline_stages_2_WAYS_TAGS_2_fault <= load_pipeline_stages_1_WAYS_TAGS_2_fault;
    load_pipeline_stages_2_WAYS_TAGS_3_loaded <= load_pipeline_stages_1_WAYS_TAGS_3_loaded;
    load_pipeline_stages_2_WAYS_TAGS_3_address <= load_pipeline_stages_1_WAYS_TAGS_3_address;
    load_pipeline_stages_2_WAYS_TAGS_3_fault <= load_pipeline_stages_1_WAYS_TAGS_3_fault;
    load_pipeline_stages_2_WAYS_HITS <= load_pipeline_stages_1_WAYS_HITS;
    load_pipeline_stages_2_STATUS_0_dirty <= load_pipeline_stages_1_STATUS_overloaded_0_dirty;
    load_pipeline_stages_2_STATUS_1_dirty <= load_pipeline_stages_1_STATUS_overloaded_1_dirty;
    load_pipeline_stages_2_STATUS_2_dirty <= load_pipeline_stages_1_STATUS_overloaded_2_dirty;
    load_pipeline_stages_2_STATUS_3_dirty <= load_pipeline_stages_1_STATUS_overloaded_3_dirty;
    load_pipeline_stages_2_LOCKED <= load_pipeline_stages_1_LOCKED;
    load_pipeline_stages_2_NEED_UNIQUE <= load_pipeline_stages_1_NEED_UNIQUE;
    store_pipeline_stages_1_ADDRESS_POST_TRANSLATION <= store_pipeline_stages_0_ADDRESS_POST_TRANSLATION;
    store_pipeline_stages_1_CPU_WORD <= store_pipeline_stages_0_CPU_WORD;
    store_pipeline_stages_1_CPU_MASK <= store_pipeline_stages_0_CPU_MASK;
    store_pipeline_stages_1_IO <= store_pipeline_stages_0_IO;
    store_pipeline_stages_1_FLUSH <= store_pipeline_stages_0_FLUSH;
    store_pipeline_stages_1_FLUSH_FREE <= store_pipeline_stages_0_FLUSH_FREE;
    store_pipeline_stages_1_PREFETCH <= store_pipeline_stages_0_PREFETCH;
    store_pipeline_stages_1_GENERATION <= store_pipeline_stages_0_GENERATION;
    store_pipeline_stages_1_WAYS_HAZARD <= store_pipeline_stages_0_WAYS_HAZARD;
    store_pipeline_stages_2_WAYS_HAZARD <= store_pipeline_stages_1_WAYS_HAZARD_overloaded;
    store_pipeline_stages_2_ADDRESS_POST_TRANSLATION <= store_pipeline_stages_1_ADDRESS_POST_TRANSLATION;
    store_pipeline_stages_2_PLRU_0 <= store_pipeline_stages_1_PLRU_0;
    store_pipeline_stages_2_PLRU_1 <= store_pipeline_stages_1_PLRU_1;
    store_pipeline_stages_2_WAYS_TAGS_0_loaded <= store_pipeline_stages_1_WAYS_TAGS_0_loaded;
    store_pipeline_stages_2_WAYS_TAGS_0_address <= store_pipeline_stages_1_WAYS_TAGS_0_address;
    store_pipeline_stages_2_WAYS_TAGS_0_fault <= store_pipeline_stages_1_WAYS_TAGS_0_fault;
    store_pipeline_stages_2_WAYS_TAGS_1_loaded <= store_pipeline_stages_1_WAYS_TAGS_1_loaded;
    store_pipeline_stages_2_WAYS_TAGS_1_address <= store_pipeline_stages_1_WAYS_TAGS_1_address;
    store_pipeline_stages_2_WAYS_TAGS_1_fault <= store_pipeline_stages_1_WAYS_TAGS_1_fault;
    store_pipeline_stages_2_WAYS_TAGS_2_loaded <= store_pipeline_stages_1_WAYS_TAGS_2_loaded;
    store_pipeline_stages_2_WAYS_TAGS_2_address <= store_pipeline_stages_1_WAYS_TAGS_2_address;
    store_pipeline_stages_2_WAYS_TAGS_2_fault <= store_pipeline_stages_1_WAYS_TAGS_2_fault;
    store_pipeline_stages_2_WAYS_TAGS_3_loaded <= store_pipeline_stages_1_WAYS_TAGS_3_loaded;
    store_pipeline_stages_2_WAYS_TAGS_3_address <= store_pipeline_stages_1_WAYS_TAGS_3_address;
    store_pipeline_stages_2_WAYS_TAGS_3_fault <= store_pipeline_stages_1_WAYS_TAGS_3_fault;
    store_pipeline_stages_2_WAYS_HITS <= store_pipeline_stages_1_WAYS_HITS;
    store_pipeline_stages_2_WAYS_HIT <= store_pipeline_stages_1_WAYS_HIT;
    store_pipeline_stages_2_STATUS_0_dirty <= store_pipeline_stages_1_STATUS_overloaded_0_dirty;
    store_pipeline_stages_2_STATUS_1_dirty <= store_pipeline_stages_1_STATUS_overloaded_1_dirty;
    store_pipeline_stages_2_STATUS_2_dirty <= store_pipeline_stages_1_STATUS_overloaded_2_dirty;
    store_pipeline_stages_2_STATUS_3_dirty <= store_pipeline_stages_1_STATUS_overloaded_3_dirty;
    store_pipeline_stages_2_REFILL_HITS_EARLY <= store_pipeline_stages_1_REFILL_HITS_EARLY;
    store_pipeline_stages_2_GENERATION <= store_pipeline_stages_1_GENERATION;
    store_pipeline_stages_2_PREFETCH <= store_pipeline_stages_1_PREFETCH;
    store_pipeline_stages_2_FLUSH <= store_pipeline_stages_1_FLUSH;
    store_pipeline_stages_2_IO <= store_pipeline_stages_1_IO;
    store_pipeline_stages_2_CPU_WORD <= store_pipeline_stages_1_CPU_WORD;
    store_pipeline_stages_2_CPU_MASK <= store_pipeline_stages_1_CPU_MASK;
    store_pipeline_stages_2_FLUSH_FREE <= store_pipeline_stages_1_FLUSH_FREE;
    if(banks_0_read_cmd_valid) begin
      _zz_39 <= banks_0_write_payload_mask;
    end
    if(banks_1_read_cmd_valid) begin
      _zz_40 <= banks_1_write_payload_mask;
    end
    if(banks_2_read_cmd_valid) begin
      _zz_41 <= banks_2_write_payload_mask;
    end
    if(banks_3_read_cmd_valid) begin
      _zz_42 <= banks_3_write_payload_mask;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      status_writeLast_valid <= 1'b0;
      wayRandom_value <= 2'b00;
      invalidate_counter <= 7'h00;
      invalidate_firstEver <= 1'b1;
      refill_slots_0_valid <= 1'b0;
      refill_slots_1_valid <= 1'b0;
      refill_pushCounter <= 32'h00000000;
      refill_read_arbiter_lock <= 2'b00;
      refill_read_wordIndex <= 3'b000;
      refill_read_hadError <= 1'b0;
      writeback_slots_0_valid <= 1'b0;
      writeback_slots_1_valid <= 1'b0;
      writeback_read_arbiter_lock <= 2'b00;
      writeback_read_wordIndex <= 3'b000;
      writeback_read_slotReadLast_valid <= 1'b0;
      writeback_write_arbiter_lock <= 2'b00;
      writeback_write_wordIndex <= 3'b000;
      writeback_write_bufferRead_rValid <= 1'b0;
      load_pipeline_stages_1_valid <= 1'b0;
      load_pipeline_stages_2_valid <= 1'b0;
      store_target <= 1'b0;
      store_pipeline_stages_1_valid <= 1'b0;
      store_pipeline_stages_2_valid <= 1'b0;
      when_MultiportRam_l328 <= 1'b0;
      when_MultiportRam_l328_1 <= 1'b0;
      when_MultiportRam_l328_2 <= 1'b0;
      when_MultiportRam_l328_3 <= 1'b0;
      when_MultiportRam_l328_4 <= 1'b0;
    end else begin
      status_writeLast_valid <= status_write_valid;
      wayRandom_value <= wayRandom_valueNext;
      if(when_DataCache_l887) begin
        invalidate_counter <= (invalidate_counter + 7'h01);
      end
      if(invalidate_done) begin
        invalidate_firstEver <= 1'b0;
      end
      if(when_DataCache_l933) begin
        refill_slots_0_valid <= 1'b0;
      end
      if(when_DataCache_l933_1) begin
        refill_slots_1_valid <= 1'b0;
      end
      if(refill_push_valid) begin
        refill_pushCounter <= (refill_pushCounter + 32'h00000001);
      end
      if(refill_push_valid) begin
        if(when_DataCache_l960) begin
          refill_slots_0_valid <= 1'b1;
        end
      end
      if(refill_push_valid) begin
        if(when_DataCache_l960_1) begin
          refill_slots_1_valid <= 1'b1;
        end
      end
      refill_read_arbiter_lock <= refill_read_arbiter_oh;
      if(when_DataCache_l985) begin
        refill_read_arbiter_lock <= 2'b00;
      end
      if(when_DataCache_l1025) begin
        refill_read_hadError <= 1'b1;
      end
      if(io_mem_read_rsp_valid) begin
        if(refill_read_rspWithData) begin
          refill_read_wordIndex <= (refill_read_wordIndex + 3'b001);
        end
        if(when_DataCache_l1036) begin
          refill_read_hadError <= 1'b0;
        end
      end
      if(writeback_slots_0_fire) begin
        writeback_slots_0_valid <= 1'b0;
      end
      if(writeback_slots_1_fire) begin
        writeback_slots_1_valid <= 1'b0;
      end
      if(writeback_push_valid) begin
        if(when_DataCache_l1127) begin
          writeback_slots_0_valid <= 1'b1;
        end
      end
      if(writeback_push_valid) begin
        if(when_DataCache_l1127_1) begin
          writeback_slots_1_valid <= 1'b1;
        end
      end
      writeback_read_arbiter_lock <= writeback_read_arbiter_oh;
      writeback_read_wordIndex <= (writeback_read_wordIndex + _zz_writeback_read_wordIndex);
      if(when_DataCache_l1174) begin
        writeback_read_arbiter_lock <= 2'b00;
      end
      writeback_read_slotReadLast_valid <= writeback_read_slotRead_valid;
      writeback_write_arbiter_lock <= writeback_write_arbiter_oh;
      writeback_write_wordIndex <= (writeback_write_wordIndex + _zz_writeback_write_wordIndex);
      if(when_DataCache_l1252) begin
        writeback_write_arbiter_lock <= 2'b00;
      end
      if(writeback_write_bufferRead_ready) begin
        writeback_write_bufferRead_rValid <= writeback_write_bufferRead_valid;
      end
      load_pipeline_stages_1_valid <= _zz_load_pipeline_stages_1_valid;
      load_pipeline_stages_2_valid <= _zz_load_pipeline_stages_2_valid;
      if(when_DataCache_l1804) begin
        store_target <= (! store_target);
      end
      store_pipeline_stages_1_valid <= _zz_store_pipeline_stages_1_valid;
      store_pipeline_stages_2_valid <= _zz_store_pipeline_stages_2_valid;
      if(banks_0_read_cmd_valid) begin
        when_MultiportRam_l328 <= (banks_0_write_valid && (banks_0_write_payload_address == banks_0_read_cmd_payload));
      end
      if(banks_1_read_cmd_valid) begin
        when_MultiportRam_l328_1 <= (banks_1_write_valid && (banks_1_write_payload_address == banks_1_read_cmd_payload));
      end
      if(banks_2_read_cmd_valid) begin
        when_MultiportRam_l328_2 <= (banks_2_write_valid && (banks_2_write_payload_address == banks_2_read_cmd_payload));
      end
      if(banks_3_read_cmd_valid) begin
        when_MultiportRam_l328_3 <= (banks_3_write_valid && (banks_3_write_payload_address == banks_3_read_cmd_payload));
      end
      if(writeback_write_bufferRead_ready) begin
        when_MultiportRam_l328_4 <= (_zz_when_MultiportRam_l328 && (_zz_when_MultiportRam_l328_1 == _zz_when_MultiportRam_l328_2));
      end
    end
  end


endmodule

module AllocatorMultiPortMem (
  input  wire          io_push_0_valid /* verilator public */ ,
  input  wire [5:0]    io_push_0_payload /* verilator public */ ,
  input  wire          io_push_1_valid /* verilator public */ ,
  input  wire [5:0]    io_push_1_payload /* verilator public */ ,
  input  wire [1:0]    io_pop_mask /* verilator public */ ,
  output wire          io_pop_ready /* verilator public */ ,
  input  wire          io_pop_fire /* verilator public */ ,
  output wire [5:0]    io_pop_values_0 /* verilator public */ ,
  output wire [5:0]    io_pop_values_1 /* verilator public */ ,
  input  wire          clk,
  input  wire          reset
);

  wire       [5:0]    _zz_ways_0_mem_port1;
  wire       [5:0]    _zz_ways_1_mem_port1;
  reg        [1:0]    _zz_popMaskCount;
  wire       [1:0]    _zz_popMaskCount_1;
  reg        [1:0]    _zz_ptr_pushCount;
  wire       [1:0]    _zz_ptr_pushCount_1;
  wire       [6:0]    _zz_ptr_push;
  wire       [6:0]    _zz_ptr_pop;
  wire       [6:0]    _zz_ptr_occupancy;
  wire       [6:0]    _zz_ptr_occupancy_1;
  wire       [6:0]    _zz_ptr_occupancy_2;
  wire       [1:0]    _zz_ptr_occupancy_3;
  wire       [6:0]    _zz_pushArbitration_pushOffset_1;
  wire       [0:0]    _zz_pushArbitration_pushOffset_1_1;
  wire       [6:0]    _zz_pushArbitration_pushOffset_2;
  wire       [0:0]    _zz_pushArbitration_pushOffset_2_1;
  wire       [4:0]    _zz_ways_0_mem_port;
  wire       [5:0]    _zz_ways_0_mem_port_1;
  wire                _zz_ways_0_mem_port_2;
  wire       [4:0]    _zz_ways_1_mem_port;
  wire       [5:0]    _zz_ways_1_mem_port_1;
  wire                _zz_ways_1_mem_port_2;
  reg        [5:0]    _zz_io_pop_values_0;
  wire       [0:0]    _zz_io_pop_values_0_1;
  wire       [6:0]    _zz_popArbitration_popOffset_1;
  wire       [0:0]    _zz_popArbitration_popOffset_1_1;
  reg        [5:0]    _zz_io_pop_values_1;
  wire       [0:0]    _zz_io_pop_values_1_1;
  wire       [6:0]    _zz_popArbitration_popOffset_2;
  wire       [0:0]    _zz_popArbitration_popOffset_2_1;
  reg        [6:0]    popArbitration_popOffset_2;
  reg        [6:0]    popArbitration_popOffset_1;
  reg        [6:0]    pushArbitration_pushOffset_2;
  reg        [6:0]    pushArbitration_pushOffset_1;
  wire       [1:0]    popMaskCount;
  reg        [6:0]    ptr_push;
  reg        [6:0]    ptr_pop;
  reg        [6:0]    ptr_occupancy;
  wire       [1:0]    ptr_pushCount;
  wire       [6:0]    pushArbitration_pushOffset;
  wire       [6:0]    pushArbitration_push_0_ptr;
  wire       [6:0]    pushArbitration_push_1_ptr;
  wire       [6:0]    ways_0_push_offset;
  wire       [1:0]    ways_0_push_hits;
  wire       [6:0]    ways_0_pop_offset;
  wire       [4:0]    _zz_ways_0_pop_data;
  wire       [5:0]    ways_0_pop_data;
  wire       [6:0]    ways_1_push_offset;
  wire       [1:0]    ways_1_push_hits;
  wire       [6:0]    ways_1_pop_offset;
  wire       [4:0]    _zz_ways_1_pop_data;
  wire       [5:0]    ways_1_pop_data;
  wire       [6:0]    popArbitration_popOffset;
  wire       [6:0]    popArbitration_pop_0_ptr;
  wire       [6:0]    popArbitration_pop_1_ptr;
  (* ram_style = "distributed" *) reg [5:0] ways_0_mem [0:31];
  (* ram_style = "distributed" *) reg [5:0] ways_1_mem [0:31];

  assign _zz_ptr_push = {5'd0, ptr_pushCount};
  assign _zz_ptr_pop = {5'd0, popMaskCount};
  assign _zz_ptr_occupancy = (ptr_occupancy + _zz_ptr_occupancy_1);
  assign _zz_ptr_occupancy_1 = {5'd0, ptr_pushCount};
  assign _zz_ptr_occupancy_3 = (io_pop_fire ? popMaskCount : 2'b00);
  assign _zz_ptr_occupancy_2 = {5'd0, _zz_ptr_occupancy_3};
  assign _zz_pushArbitration_pushOffset_1_1 = io_push_0_valid;
  assign _zz_pushArbitration_pushOffset_1 = {6'd0, _zz_pushArbitration_pushOffset_1_1};
  assign _zz_pushArbitration_pushOffset_2_1 = io_push_1_valid;
  assign _zz_pushArbitration_pushOffset_2 = {6'd0, _zz_pushArbitration_pushOffset_2_1};
  assign _zz_popArbitration_popOffset_1_1 = io_pop_mask[0];
  assign _zz_popArbitration_popOffset_1 = {6'd0, _zz_popArbitration_popOffset_1_1};
  assign _zz_popArbitration_popOffset_2_1 = io_pop_mask[1];
  assign _zz_popArbitration_popOffset_2 = {6'd0, _zz_popArbitration_popOffset_2_1};
  assign _zz_ways_0_mem_port = ways_0_push_offset[5 : 1];
  assign _zz_ways_0_mem_port_1 = (ways_0_push_hits[0] ? io_push_0_payload : io_push_1_payload);
  assign _zz_ways_0_mem_port_2 = (|ways_0_push_hits);
  assign _zz_ways_1_mem_port = ways_1_push_offset[5 : 1];
  assign _zz_ways_1_mem_port_1 = (ways_1_push_hits[0] ? io_push_0_payload : io_push_1_payload);
  assign _zz_ways_1_mem_port_2 = (|ways_1_push_hits);
  assign _zz_popMaskCount_1 = {io_pop_mask[1],io_pop_mask[0]};
  assign _zz_ptr_pushCount_1 = {io_push_1_valid,io_push_0_valid};
  assign _zz_io_pop_values_0_1 = popArbitration_pop_0_ptr[0 : 0];
  assign _zz_io_pop_values_1_1 = popArbitration_pop_1_ptr[0 : 0];
  always @(posedge clk) begin
    if(_zz_ways_0_mem_port_2) begin
      ways_0_mem[_zz_ways_0_mem_port] <= _zz_ways_0_mem_port_1;
    end
  end

  assign _zz_ways_0_mem_port1 = ways_0_mem[_zz_ways_0_pop_data];
  always @(posedge clk) begin
    if(_zz_ways_1_mem_port_2) begin
      ways_1_mem[_zz_ways_1_mem_port] <= _zz_ways_1_mem_port_1;
    end
  end

  assign _zz_ways_1_mem_port1 = ways_1_mem[_zz_ways_1_pop_data];
  always @(*) begin
    case(_zz_popMaskCount_1)
      2'b00 : _zz_popMaskCount = 2'b00;
      2'b01 : _zz_popMaskCount = 2'b01;
      2'b10 : _zz_popMaskCount = 2'b01;
      default : _zz_popMaskCount = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_ptr_pushCount_1)
      2'b00 : _zz_ptr_pushCount = 2'b00;
      2'b01 : _zz_ptr_pushCount = 2'b01;
      2'b10 : _zz_ptr_pushCount = 2'b01;
      default : _zz_ptr_pushCount = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_io_pop_values_0_1)
      1'b0 : _zz_io_pop_values_0 = ways_0_pop_data;
      default : _zz_io_pop_values_0 = ways_1_pop_data;
    endcase
  end

  always @(*) begin
    case(_zz_io_pop_values_1_1)
      1'b0 : _zz_io_pop_values_1 = ways_0_pop_data;
      default : _zz_io_pop_values_1 = ways_1_pop_data;
    endcase
  end

  always @(*) begin
    popArbitration_popOffset_2 = popArbitration_popOffset_1;
    popArbitration_popOffset_2 = (popArbitration_popOffset_1 + _zz_popArbitration_popOffset_2);
  end

  always @(*) begin
    popArbitration_popOffset_1 = popArbitration_popOffset;
    popArbitration_popOffset_1 = (popArbitration_popOffset + _zz_popArbitration_popOffset_1);
  end

  always @(*) begin
    pushArbitration_pushOffset_2 = pushArbitration_pushOffset_1;
    pushArbitration_pushOffset_2 = (pushArbitration_pushOffset_1 + _zz_pushArbitration_pushOffset_2);
  end

  always @(*) begin
    pushArbitration_pushOffset_1 = pushArbitration_pushOffset;
    pushArbitration_pushOffset_1 = (pushArbitration_pushOffset + _zz_pushArbitration_pushOffset_1);
  end

  assign popMaskCount = _zz_popMaskCount;
  assign ptr_pushCount = _zz_ptr_pushCount;
  assign pushArbitration_pushOffset = ptr_push;
  assign pushArbitration_push_0_ptr = pushArbitration_pushOffset;
  assign pushArbitration_push_1_ptr = pushArbitration_pushOffset_1;
  assign ways_0_push_offset = (ptr_push + 7'h01);
  assign ways_0_push_hits = ({io_push_1_valid,io_push_0_valid} & {(pushArbitration_push_1_ptr[0 : 0] == 1'b0),(pushArbitration_push_0_ptr[0 : 0] == 1'b0)});
  assign ways_0_pop_offset = (ptr_pop + 7'h01);
  assign _zz_ways_0_pop_data = ways_0_pop_offset[5 : 1];
  assign ways_0_pop_data = _zz_ways_0_mem_port1;
  assign ways_1_push_offset = (ptr_push + 7'h00);
  assign ways_1_push_hits = ({io_push_1_valid,io_push_0_valid} & {(pushArbitration_push_1_ptr[0 : 0] == 1'b1),(pushArbitration_push_0_ptr[0 : 0] == 1'b1)});
  assign ways_1_pop_offset = (ptr_pop + 7'h00);
  assign _zz_ways_1_pop_data = ways_1_pop_offset[5 : 1];
  assign ways_1_pop_data = _zz_ways_1_mem_port1;
  assign popArbitration_popOffset = ptr_pop;
  assign popArbitration_pop_0_ptr = popArbitration_popOffset;
  assign io_pop_values_0 = _zz_io_pop_values_0;
  assign popArbitration_pop_1_ptr = popArbitration_popOffset_1;
  assign io_pop_values_1 = _zz_io_pop_values_1;
  assign io_pop_ready = (7'h02 <= ptr_occupancy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      ptr_push <= 7'h00;
      ptr_pop <= 7'h00;
      ptr_occupancy <= 7'h00;
    end else begin
      ptr_push <= (ptr_push + _zz_ptr_push);
      if(io_pop_fire) begin
        ptr_pop <= (ptr_pop + _zz_ptr_pop);
      end
      ptr_occupancy <= (_zz_ptr_occupancy - _zz_ptr_occupancy_2);
    end
  end


endmodule

module TranslatorWithRollback (
  input  wire          io_rollback,
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_payload_address,
  input  wire [5:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [4:0]    io_writes_1_payload_address,
  input  wire [5:0]    io_writes_1_payload_data,
  input  wire          io_commits_0_valid,
  input  wire [4:0]    io_commits_0_payload_address,
  input  wire [5:0]    io_commits_0_payload_data,
  input  wire          io_commits_1_valid,
  input  wire [4:0]    io_commits_1_payload_address,
  input  wire [5:0]    io_commits_1_payload_data,
  input  wire          io_reads_0_cmd_valid,
  input  wire [4:0]    io_reads_0_cmd_payload,
  output wire          io_reads_0_rsp_valid,
  output wire [5:0]    io_reads_0_rsp_payload,
  input  wire          io_reads_1_cmd_valid,
  input  wire [4:0]    io_reads_1_cmd_payload,
  output wire          io_reads_1_rsp_valid,
  output wire [5:0]    io_reads_1_rsp_payload,
  input  wire          io_reads_2_cmd_valid,
  input  wire [4:0]    io_reads_2_cmd_payload,
  output wire          io_reads_2_rsp_valid,
  output wire [5:0]    io_reads_2_rsp_payload,
  input  wire          io_reads_3_cmd_valid,
  input  wire [4:0]    io_reads_3_cmd_payload,
  output wire          io_reads_3_rsp_valid,
  output wire [5:0]    io_reads_3_rsp_payload,
  input  wire          io_reads_4_cmd_valid,
  input  wire [4:0]    io_reads_4_cmd_payload,
  output wire          io_reads_4_rsp_valid,
  output wire [5:0]    io_reads_4_rsp_payload,
  input  wire          io_reads_5_cmd_valid,
  input  wire [4:0]    io_reads_5_cmd_payload,
  output wire          io_reads_5_rsp_valid,
  output wire [5:0]    io_reads_5_rsp_payload,
  input  wire          clk,
  input  wire          reset
);

  wire                writes_ram_io_writes_0_valid;
  wire       [5:0]    writes_ram_io_writes_0_payload_data;
  wire                writes_ram_io_writes_1_valid;
  wire       [5:0]    writes_ram_io_writes_1_payload_data;
  wire                writes_ram_io_read_0_cmd_valid;
  wire                writes_ram_io_read_1_cmd_valid;
  wire                writes_ram_io_read_2_cmd_valid;
  wire                writes_ram_io_read_3_cmd_valid;
  wire                writes_ram_io_read_4_cmd_valid;
  wire                writes_ram_io_read_5_cmd_valid;
  wire                commits_ram_io_writes_0_valid;
  wire       [5:0]    commits_ram_io_writes_0_payload_data;
  wire                commits_ram_io_writes_1_valid;
  wire       [5:0]    commits_ram_io_writes_1_payload_data;
  wire                commits_ram_io_read_0_cmd_valid;
  wire                commits_ram_io_read_1_cmd_valid;
  wire                commits_ram_io_read_2_cmd_valid;
  wire                commits_ram_io_read_3_cmd_valid;
  wire                commits_ram_io_read_4_cmd_valid;
  wire                commits_ram_io_read_5_cmd_valid;
  wire       [5:0]    writes_ram_io_read_0_rsp;
  wire       [5:0]    writes_ram_io_read_1_rsp;
  wire       [5:0]    writes_ram_io_read_2_rsp;
  wire       [5:0]    writes_ram_io_read_3_rsp;
  wire       [5:0]    writes_ram_io_read_4_rsp;
  wire       [5:0]    writes_ram_io_read_5_rsp;
  wire       [5:0]    commits_ram_io_read_0_rsp;
  wire       [5:0]    commits_ram_io_read_1_rsp;
  wire       [5:0]    commits_ram_io_read_2_rsp;
  wire       [5:0]    commits_ram_io_read_3_rsp;
  wire       [5:0]    commits_ram_io_read_4_rsp;
  wire       [5:0]    commits_ram_io_read_5_rsp;
  reg        [31:0]   location_updated;
  wire                location_set_0_hits_0;
  wire                location_set_0_hits_1;
  wire                when_RfTranslationPlugin_l71;
  wire                location_set_1_hits_0;
  wire                location_set_1_hits_1;
  wire                when_RfTranslationPlugin_l71_1;
  wire                location_set_2_hits_0;
  wire                location_set_2_hits_1;
  wire                when_RfTranslationPlugin_l71_2;
  wire                location_set_3_hits_0;
  wire                location_set_3_hits_1;
  wire                when_RfTranslationPlugin_l71_3;
  wire                location_set_4_hits_0;
  wire                location_set_4_hits_1;
  wire                when_RfTranslationPlugin_l71_4;
  wire                location_set_5_hits_0;
  wire                location_set_5_hits_1;
  wire                when_RfTranslationPlugin_l71_5;
  wire                location_set_6_hits_0;
  wire                location_set_6_hits_1;
  wire                when_RfTranslationPlugin_l71_6;
  wire                location_set_7_hits_0;
  wire                location_set_7_hits_1;
  wire                when_RfTranslationPlugin_l71_7;
  wire                location_set_8_hits_0;
  wire                location_set_8_hits_1;
  wire                when_RfTranslationPlugin_l71_8;
  wire                location_set_9_hits_0;
  wire                location_set_9_hits_1;
  wire                when_RfTranslationPlugin_l71_9;
  wire                location_set_10_hits_0;
  wire                location_set_10_hits_1;
  wire                when_RfTranslationPlugin_l71_10;
  wire                location_set_11_hits_0;
  wire                location_set_11_hits_1;
  wire                when_RfTranslationPlugin_l71_11;
  wire                location_set_12_hits_0;
  wire                location_set_12_hits_1;
  wire                when_RfTranslationPlugin_l71_12;
  wire                location_set_13_hits_0;
  wire                location_set_13_hits_1;
  wire                when_RfTranslationPlugin_l71_13;
  wire                location_set_14_hits_0;
  wire                location_set_14_hits_1;
  wire                when_RfTranslationPlugin_l71_14;
  wire                location_set_15_hits_0;
  wire                location_set_15_hits_1;
  wire                when_RfTranslationPlugin_l71_15;
  wire                location_set_16_hits_0;
  wire                location_set_16_hits_1;
  wire                when_RfTranslationPlugin_l71_16;
  wire                location_set_17_hits_0;
  wire                location_set_17_hits_1;
  wire                when_RfTranslationPlugin_l71_17;
  wire                location_set_18_hits_0;
  wire                location_set_18_hits_1;
  wire                when_RfTranslationPlugin_l71_18;
  wire                location_set_19_hits_0;
  wire                location_set_19_hits_1;
  wire                when_RfTranslationPlugin_l71_19;
  wire                location_set_20_hits_0;
  wire                location_set_20_hits_1;
  wire                when_RfTranslationPlugin_l71_20;
  wire                location_set_21_hits_0;
  wire                location_set_21_hits_1;
  wire                when_RfTranslationPlugin_l71_21;
  wire                location_set_22_hits_0;
  wire                location_set_22_hits_1;
  wire                when_RfTranslationPlugin_l71_22;
  wire                location_set_23_hits_0;
  wire                location_set_23_hits_1;
  wire                when_RfTranslationPlugin_l71_23;
  wire                location_set_24_hits_0;
  wire                location_set_24_hits_1;
  wire                when_RfTranslationPlugin_l71_24;
  wire                location_set_25_hits_0;
  wire                location_set_25_hits_1;
  wire                when_RfTranslationPlugin_l71_25;
  wire                location_set_26_hits_0;
  wire                location_set_26_hits_1;
  wire                when_RfTranslationPlugin_l71_26;
  wire                location_set_27_hits_0;
  wire                location_set_27_hits_1;
  wire                when_RfTranslationPlugin_l71_27;
  wire                location_set_28_hits_0;
  wire                location_set_28_hits_1;
  wire                when_RfTranslationPlugin_l71_28;
  wire                location_set_29_hits_0;
  wire                location_set_29_hits_1;
  wire                when_RfTranslationPlugin_l71_29;
  wire                location_set_30_hits_0;
  wire                location_set_30_hits_1;
  wire                when_RfTranslationPlugin_l71_30;
  wire                location_set_31_hits_0;
  wire                location_set_31_hits_1;
  wire                when_RfTranslationPlugin_l71_31;
  wire       [5:0]    read_0_written;
  wire       [5:0]    read_0_commited;
  wire                read_0_sel;
  wire       [5:0]    read_0_muxed;
  wire       [5:0]    read_1_written;
  wire       [5:0]    read_1_commited;
  wire                read_1_sel;
  wire       [5:0]    read_1_muxed;
  wire       [5:0]    read_2_written;
  wire       [5:0]    read_2_commited;
  wire                read_2_sel;
  wire       [5:0]    read_2_muxed;
  wire       [5:0]    read_3_written;
  wire       [5:0]    read_3_commited;
  wire                read_3_sel;
  wire       [5:0]    read_3_muxed;
  wire       [5:0]    read_4_written;
  wire       [5:0]    read_4_commited;
  wire                read_4_sel;
  wire       [5:0]    read_4_muxed;
  wire       [5:0]    read_5_written;
  wire       [5:0]    read_5_commited;
  wire                read_5_sel;
  wire       [5:0]    read_5_muxed;

  RamAsyncMwXor_13 writes_ram (
    .io_writes_0_valid           (writes_ram_io_writes_0_valid            ), //i
    .io_writes_0_payload_address (io_writes_0_payload_address[4:0]        ), //i
    .io_writes_0_payload_data    (writes_ram_io_writes_0_payload_data[5:0]), //i
    .io_writes_1_valid           (writes_ram_io_writes_1_valid            ), //i
    .io_writes_1_payload_address (io_writes_1_payload_address[4:0]        ), //i
    .io_writes_1_payload_data    (writes_ram_io_writes_1_payload_data[5:0]), //i
    .io_read_0_cmd_valid         (writes_ram_io_read_0_cmd_valid          ), //i
    .io_read_0_cmd_payload       (io_reads_0_cmd_payload[4:0]             ), //i
    .io_read_0_rsp               (writes_ram_io_read_0_rsp[5:0]           ), //o
    .io_read_1_cmd_valid         (writes_ram_io_read_1_cmd_valid          ), //i
    .io_read_1_cmd_payload       (io_reads_1_cmd_payload[4:0]             ), //i
    .io_read_1_rsp               (writes_ram_io_read_1_rsp[5:0]           ), //o
    .io_read_2_cmd_valid         (writes_ram_io_read_2_cmd_valid          ), //i
    .io_read_2_cmd_payload       (io_reads_2_cmd_payload[4:0]             ), //i
    .io_read_2_rsp               (writes_ram_io_read_2_rsp[5:0]           ), //o
    .io_read_3_cmd_valid         (writes_ram_io_read_3_cmd_valid          ), //i
    .io_read_3_cmd_payload       (io_reads_3_cmd_payload[4:0]             ), //i
    .io_read_3_rsp               (writes_ram_io_read_3_rsp[5:0]           ), //o
    .io_read_4_cmd_valid         (writes_ram_io_read_4_cmd_valid          ), //i
    .io_read_4_cmd_payload       (io_reads_4_cmd_payload[4:0]             ), //i
    .io_read_4_rsp               (writes_ram_io_read_4_rsp[5:0]           ), //o
    .io_read_5_cmd_valid         (writes_ram_io_read_5_cmd_valid          ), //i
    .io_read_5_cmd_payload       (io_reads_5_cmd_payload[4:0]             ), //i
    .io_read_5_rsp               (writes_ram_io_read_5_rsp[5:0]           ), //o
    .clk                         (clk                                     ), //i
    .reset                       (reset                                   )  //i
  );
  RamAsyncMwXor_13 commits_ram (
    .io_writes_0_valid           (commits_ram_io_writes_0_valid            ), //i
    .io_writes_0_payload_address (io_commits_0_payload_address[4:0]        ), //i
    .io_writes_0_payload_data    (commits_ram_io_writes_0_payload_data[5:0]), //i
    .io_writes_1_valid           (commits_ram_io_writes_1_valid            ), //i
    .io_writes_1_payload_address (io_commits_1_payload_address[4:0]        ), //i
    .io_writes_1_payload_data    (commits_ram_io_writes_1_payload_data[5:0]), //i
    .io_read_0_cmd_valid         (commits_ram_io_read_0_cmd_valid          ), //i
    .io_read_0_cmd_payload       (io_reads_0_cmd_payload[4:0]              ), //i
    .io_read_0_rsp               (commits_ram_io_read_0_rsp[5:0]           ), //o
    .io_read_1_cmd_valid         (commits_ram_io_read_1_cmd_valid          ), //i
    .io_read_1_cmd_payload       (io_reads_1_cmd_payload[4:0]              ), //i
    .io_read_1_rsp               (commits_ram_io_read_1_rsp[5:0]           ), //o
    .io_read_2_cmd_valid         (commits_ram_io_read_2_cmd_valid          ), //i
    .io_read_2_cmd_payload       (io_reads_2_cmd_payload[4:0]              ), //i
    .io_read_2_rsp               (commits_ram_io_read_2_rsp[5:0]           ), //o
    .io_read_3_cmd_valid         (commits_ram_io_read_3_cmd_valid          ), //i
    .io_read_3_cmd_payload       (io_reads_3_cmd_payload[4:0]              ), //i
    .io_read_3_rsp               (commits_ram_io_read_3_rsp[5:0]           ), //o
    .io_read_4_cmd_valid         (commits_ram_io_read_4_cmd_valid          ), //i
    .io_read_4_cmd_payload       (io_reads_4_cmd_payload[4:0]              ), //i
    .io_read_4_rsp               (commits_ram_io_read_4_rsp[5:0]           ), //o
    .io_read_5_cmd_valid         (commits_ram_io_read_5_cmd_valid          ), //i
    .io_read_5_cmd_payload       (io_reads_5_cmd_payload[4:0]              ), //i
    .io_read_5_rsp               (commits_ram_io_read_5_rsp[5:0]           ), //o
    .clk                         (clk                                      ), //i
    .reset                       (reset                                    )  //i
  );
  assign location_set_0_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h00));
  assign location_set_0_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h00));
  assign when_RfTranslationPlugin_l71 = ({location_set_0_hits_1,location_set_0_hits_0} != 2'b00);
  assign location_set_1_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h01));
  assign location_set_1_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h01));
  assign when_RfTranslationPlugin_l71_1 = ({location_set_1_hits_1,location_set_1_hits_0} != 2'b00);
  assign location_set_2_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h02));
  assign location_set_2_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h02));
  assign when_RfTranslationPlugin_l71_2 = ({location_set_2_hits_1,location_set_2_hits_0} != 2'b00);
  assign location_set_3_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h03));
  assign location_set_3_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h03));
  assign when_RfTranslationPlugin_l71_3 = ({location_set_3_hits_1,location_set_3_hits_0} != 2'b00);
  assign location_set_4_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h04));
  assign location_set_4_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h04));
  assign when_RfTranslationPlugin_l71_4 = ({location_set_4_hits_1,location_set_4_hits_0} != 2'b00);
  assign location_set_5_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h05));
  assign location_set_5_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h05));
  assign when_RfTranslationPlugin_l71_5 = ({location_set_5_hits_1,location_set_5_hits_0} != 2'b00);
  assign location_set_6_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h06));
  assign location_set_6_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h06));
  assign when_RfTranslationPlugin_l71_6 = ({location_set_6_hits_1,location_set_6_hits_0} != 2'b00);
  assign location_set_7_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h07));
  assign location_set_7_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h07));
  assign when_RfTranslationPlugin_l71_7 = ({location_set_7_hits_1,location_set_7_hits_0} != 2'b00);
  assign location_set_8_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h08));
  assign location_set_8_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h08));
  assign when_RfTranslationPlugin_l71_8 = ({location_set_8_hits_1,location_set_8_hits_0} != 2'b00);
  assign location_set_9_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h09));
  assign location_set_9_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h09));
  assign when_RfTranslationPlugin_l71_9 = ({location_set_9_hits_1,location_set_9_hits_0} != 2'b00);
  assign location_set_10_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0a));
  assign location_set_10_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h0a));
  assign when_RfTranslationPlugin_l71_10 = ({location_set_10_hits_1,location_set_10_hits_0} != 2'b00);
  assign location_set_11_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0b));
  assign location_set_11_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h0b));
  assign when_RfTranslationPlugin_l71_11 = ({location_set_11_hits_1,location_set_11_hits_0} != 2'b00);
  assign location_set_12_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0c));
  assign location_set_12_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h0c));
  assign when_RfTranslationPlugin_l71_12 = ({location_set_12_hits_1,location_set_12_hits_0} != 2'b00);
  assign location_set_13_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0d));
  assign location_set_13_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h0d));
  assign when_RfTranslationPlugin_l71_13 = ({location_set_13_hits_1,location_set_13_hits_0} != 2'b00);
  assign location_set_14_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0e));
  assign location_set_14_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h0e));
  assign when_RfTranslationPlugin_l71_14 = ({location_set_14_hits_1,location_set_14_hits_0} != 2'b00);
  assign location_set_15_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h0f));
  assign location_set_15_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h0f));
  assign when_RfTranslationPlugin_l71_15 = ({location_set_15_hits_1,location_set_15_hits_0} != 2'b00);
  assign location_set_16_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h10));
  assign location_set_16_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h10));
  assign when_RfTranslationPlugin_l71_16 = ({location_set_16_hits_1,location_set_16_hits_0} != 2'b00);
  assign location_set_17_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h11));
  assign location_set_17_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h11));
  assign when_RfTranslationPlugin_l71_17 = ({location_set_17_hits_1,location_set_17_hits_0} != 2'b00);
  assign location_set_18_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h12));
  assign location_set_18_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h12));
  assign when_RfTranslationPlugin_l71_18 = ({location_set_18_hits_1,location_set_18_hits_0} != 2'b00);
  assign location_set_19_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h13));
  assign location_set_19_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h13));
  assign when_RfTranslationPlugin_l71_19 = ({location_set_19_hits_1,location_set_19_hits_0} != 2'b00);
  assign location_set_20_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h14));
  assign location_set_20_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h14));
  assign when_RfTranslationPlugin_l71_20 = ({location_set_20_hits_1,location_set_20_hits_0} != 2'b00);
  assign location_set_21_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h15));
  assign location_set_21_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h15));
  assign when_RfTranslationPlugin_l71_21 = ({location_set_21_hits_1,location_set_21_hits_0} != 2'b00);
  assign location_set_22_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h16));
  assign location_set_22_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h16));
  assign when_RfTranslationPlugin_l71_22 = ({location_set_22_hits_1,location_set_22_hits_0} != 2'b00);
  assign location_set_23_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h17));
  assign location_set_23_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h17));
  assign when_RfTranslationPlugin_l71_23 = ({location_set_23_hits_1,location_set_23_hits_0} != 2'b00);
  assign location_set_24_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h18));
  assign location_set_24_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h18));
  assign when_RfTranslationPlugin_l71_24 = ({location_set_24_hits_1,location_set_24_hits_0} != 2'b00);
  assign location_set_25_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h19));
  assign location_set_25_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h19));
  assign when_RfTranslationPlugin_l71_25 = ({location_set_25_hits_1,location_set_25_hits_0} != 2'b00);
  assign location_set_26_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1a));
  assign location_set_26_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h1a));
  assign when_RfTranslationPlugin_l71_26 = ({location_set_26_hits_1,location_set_26_hits_0} != 2'b00);
  assign location_set_27_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1b));
  assign location_set_27_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h1b));
  assign when_RfTranslationPlugin_l71_27 = ({location_set_27_hits_1,location_set_27_hits_0} != 2'b00);
  assign location_set_28_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1c));
  assign location_set_28_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h1c));
  assign when_RfTranslationPlugin_l71_28 = ({location_set_28_hits_1,location_set_28_hits_0} != 2'b00);
  assign location_set_29_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1d));
  assign location_set_29_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h1d));
  assign when_RfTranslationPlugin_l71_29 = ({location_set_29_hits_1,location_set_29_hits_0} != 2'b00);
  assign location_set_30_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1e));
  assign location_set_30_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h1e));
  assign when_RfTranslationPlugin_l71_30 = ({location_set_30_hits_1,location_set_30_hits_0} != 2'b00);
  assign location_set_31_hits_0 = (io_writes_0_valid && (io_writes_0_payload_address == 5'h1f));
  assign location_set_31_hits_1 = (io_writes_1_valid && (io_writes_1_payload_address == 5'h1f));
  assign when_RfTranslationPlugin_l71_31 = ({location_set_31_hits_1,location_set_31_hits_0} != 2'b00);
  assign read_0_written = writes_ram_io_read_0_rsp;
  assign read_0_commited = commits_ram_io_read_0_rsp;
  assign read_0_sel = location_updated[io_reads_0_cmd_payload];
  assign read_0_muxed = (read_0_sel ? read_0_written : read_0_commited);
  assign io_reads_0_rsp_valid = io_reads_0_cmd_valid;
  assign io_reads_0_rsp_payload = read_0_muxed;
  assign read_1_written = writes_ram_io_read_1_rsp;
  assign read_1_commited = commits_ram_io_read_1_rsp;
  assign read_1_sel = location_updated[io_reads_1_cmd_payload];
  assign read_1_muxed = (read_1_sel ? read_1_written : read_1_commited);
  assign io_reads_1_rsp_valid = io_reads_1_cmd_valid;
  assign io_reads_1_rsp_payload = read_1_muxed;
  assign read_2_written = writes_ram_io_read_2_rsp;
  assign read_2_commited = commits_ram_io_read_2_rsp;
  assign read_2_sel = location_updated[io_reads_2_cmd_payload];
  assign read_2_muxed = (read_2_sel ? read_2_written : read_2_commited);
  assign io_reads_2_rsp_valid = io_reads_2_cmd_valid;
  assign io_reads_2_rsp_payload = read_2_muxed;
  assign read_3_written = writes_ram_io_read_3_rsp;
  assign read_3_commited = commits_ram_io_read_3_rsp;
  assign read_3_sel = location_updated[io_reads_3_cmd_payload];
  assign read_3_muxed = (read_3_sel ? read_3_written : read_3_commited);
  assign io_reads_3_rsp_valid = io_reads_3_cmd_valid;
  assign io_reads_3_rsp_payload = read_3_muxed;
  assign read_4_written = writes_ram_io_read_4_rsp;
  assign read_4_commited = commits_ram_io_read_4_rsp;
  assign read_4_sel = location_updated[io_reads_4_cmd_payload];
  assign read_4_muxed = (read_4_sel ? read_4_written : read_4_commited);
  assign io_reads_4_rsp_valid = io_reads_4_cmd_valid;
  assign io_reads_4_rsp_payload = read_4_muxed;
  assign read_5_written = writes_ram_io_read_5_rsp;
  assign read_5_commited = commits_ram_io_read_5_rsp;
  assign read_5_sel = location_updated[io_reads_5_cmd_payload];
  assign read_5_muxed = (read_5_sel ? read_5_written : read_5_commited);
  assign io_reads_5_rsp_valid = io_reads_5_cmd_valid;
  assign io_reads_5_rsp_payload = read_5_muxed;
  assign writes_ram_io_writes_0_valid = (io_writes_0_valid && (! ((io_writes_1_valid && (io_writes_1_payload_address == io_writes_0_payload_address)) != 1'b0)));
  assign writes_ram_io_writes_0_payload_data = io_writes_0_payload_data;
  assign writes_ram_io_writes_1_valid = (io_writes_1_valid && (! 1'b0));
  assign writes_ram_io_writes_1_payload_data = io_writes_1_payload_data;
  assign writes_ram_io_read_0_cmd_valid = 1'b1;
  assign writes_ram_io_read_1_cmd_valid = 1'b1;
  assign writes_ram_io_read_2_cmd_valid = 1'b1;
  assign writes_ram_io_read_3_cmd_valid = 1'b1;
  assign writes_ram_io_read_4_cmd_valid = 1'b1;
  assign writes_ram_io_read_5_cmd_valid = 1'b1;
  assign commits_ram_io_writes_0_valid = (io_commits_0_valid && (! ((io_commits_1_valid && (io_commits_1_payload_address == io_commits_0_payload_address)) != 1'b0)));
  assign commits_ram_io_writes_0_payload_data = io_commits_0_payload_data;
  assign commits_ram_io_writes_1_valid = (io_commits_1_valid && (! 1'b0));
  assign commits_ram_io_writes_1_payload_data = io_commits_1_payload_data;
  assign commits_ram_io_read_0_cmd_valid = 1'b1;
  assign commits_ram_io_read_1_cmd_valid = 1'b1;
  assign commits_ram_io_read_2_cmd_valid = 1'b1;
  assign commits_ram_io_read_3_cmd_valid = 1'b1;
  assign commits_ram_io_read_4_cmd_valid = 1'b1;
  assign commits_ram_io_read_5_cmd_valid = 1'b1;
  always @(posedge clk) begin
    if(when_RfTranslationPlugin_l71) begin
      location_updated[0] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_1) begin
      location_updated[1] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_2) begin
      location_updated[2] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_3) begin
      location_updated[3] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_4) begin
      location_updated[4] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_5) begin
      location_updated[5] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_6) begin
      location_updated[6] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_7) begin
      location_updated[7] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_8) begin
      location_updated[8] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_9) begin
      location_updated[9] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_10) begin
      location_updated[10] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_11) begin
      location_updated[11] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_12) begin
      location_updated[12] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_13) begin
      location_updated[13] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_14) begin
      location_updated[14] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_15) begin
      location_updated[15] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_16) begin
      location_updated[16] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_17) begin
      location_updated[17] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_18) begin
      location_updated[18] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_19) begin
      location_updated[19] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_20) begin
      location_updated[20] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_21) begin
      location_updated[21] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_22) begin
      location_updated[22] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_23) begin
      location_updated[23] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_24) begin
      location_updated[24] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_25) begin
      location_updated[25] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_26) begin
      location_updated[26] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_27) begin
      location_updated[27] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_28) begin
      location_updated[28] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_29) begin
      location_updated[29] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_30) begin
      location_updated[30] <= 1'b1;
    end
    if(when_RfTranslationPlugin_l71_31) begin
      location_updated[31] <= 1'b1;
    end
    if(io_rollback) begin
      location_updated <= 32'h00000000;
    end
  end


endmodule

//RamAsyncMwXor_8 replaced by RamAsyncMwXor_9

module RamAsyncMwXor_9 (
  input  wire          io_writes_0_valid,
  input  wire [3:0]    io_writes_0_payload_address,
  input  wire [0:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [3:0]    io_writes_1_payload_address,
  input  wire [0:0]    io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [3:0]    io_read_0_cmd_payload,
  output wire [0:0]    io_read_0_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [0:0]    _zz_ram_0_port1;
  wire       [0:0]    _zz_ram_0_port2;
  wire       [0:0]    _zz_ram_1_port0;
  wire       [0:0]    _zz_ram_1_port2;
  wire       [0:0]    writes_0_values_0;
  wire       [0:0]    writes_0_xored;
  wire       [0:0]    writes_1_values_0;
  wire       [0:0]    writes_1_xored;
  wire       [0:0]    reads_0_values_0;
  wire       [0:0]    reads_0_values_1;
  wire       [0:0]    reads_0_xored;
  (* ram_style = "distributed" *) reg [0:0] ram_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] ram_1 [0:15];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_read_0_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_xored = (io_writes_0_payload_data ^ writes_0_values_0);
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_xored = (io_writes_1_payload_data ^ writes_1_values_0);
  assign reads_0_values_0 = _zz_ram_0_port2;
  assign reads_0_values_1 = _zz_ram_1_port2;
  assign reads_0_xored = (reads_0_values_0 ^ reads_0_values_1);
  assign io_read_0_rsp = reads_0_xored;

endmodule

module RamAsyncMwXor_10 (
  input  wire          io_writes_0_valid,
  input  wire [3:0]    io_writes_0_payload_address,
  input  wire [0:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [3:0]    io_writes_1_payload_address,
  input  wire [0:0]    io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [3:0]    io_read_0_cmd_payload,
  output wire [0:0]    io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [3:0]    io_read_1_cmd_payload,
  output wire [0:0]    io_read_1_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [0:0]    _zz_ram_0_port1;
  wire       [0:0]    _zz_ram_0_port2;
  wire       [0:0]    _zz_ram_0_port3;
  wire       [0:0]    _zz_ram_1_port0;
  wire       [0:0]    _zz_ram_1_port2;
  wire       [0:0]    _zz_ram_1_port3;
  wire       [0:0]    writes_0_values_0;
  wire       [0:0]    writes_0_xored;
  wire       [0:0]    writes_1_values_0;
  wire       [0:0]    writes_1_xored;
  wire       [0:0]    reads_0_values_0;
  wire       [0:0]    reads_0_values_1;
  wire       [0:0]    reads_0_xored;
  wire       [0:0]    reads_1_values_0;
  wire       [0:0]    reads_1_values_1;
  wire       [0:0]    reads_1_xored;
  (* ram_style = "distributed" *) reg [0:0] ram_0 [0:15];
  (* ram_style = "distributed" *) reg [0:0] ram_1 [0:15];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_0_port3 = ram_0[io_read_1_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_1_port3 = ram_1[io_read_1_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_xored = (io_writes_0_payload_data ^ writes_0_values_0);
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_xored = (io_writes_1_payload_data ^ writes_1_values_0);
  assign reads_0_values_0 = _zz_ram_0_port2;
  assign reads_0_values_1 = _zz_ram_1_port2;
  assign reads_0_xored = (reads_0_values_0 ^ reads_0_values_1);
  assign io_read_0_rsp = reads_0_xored;
  assign reads_1_values_0 = _zz_ram_0_port3;
  assign reads_1_values_1 = _zz_ram_1_port3;
  assign reads_1_xored = (reads_1_values_0 ^ reads_1_values_1);
  assign io_read_1_rsp = reads_1_xored;

endmodule

module RamAsyncMwXor_12 (
  input  wire          io_writes_0_valid,
  input  wire [5:0]    io_writes_0_payload_address,
  input  wire [0:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [5:0]    io_writes_1_payload_address,
  input  wire [0:0]    io_writes_1_payload_data,
  input  wire          io_writes_2_valid,
  input  wire [5:0]    io_writes_2_payload_address,
  input  wire [0:0]    io_writes_2_payload_data,
  input  wire          io_writes_3_valid,
  input  wire [5:0]    io_writes_3_payload_address,
  input  wire [0:0]    io_writes_3_payload_data,
  input  wire          io_writes_4_valid,
  input  wire [5:0]    io_writes_4_payload_address,
  input  wire [0:0]    io_writes_4_payload_data,
  input  wire          io_writes_5_valid,
  input  wire [5:0]    io_writes_5_payload_address,
  input  wire [0:0]    io_writes_5_payload_data,
  input  wire          io_writes_6_valid,
  input  wire [5:0]    io_writes_6_payload_address,
  input  wire [0:0]    io_writes_6_payload_data,
  input  wire          io_writes_7_valid,
  input  wire [5:0]    io_writes_7_payload_address,
  input  wire [0:0]    io_writes_7_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [5:0]    io_read_0_cmd_payload,
  output wire [0:0]    io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [5:0]    io_read_1_cmd_payload,
  output wire [0:0]    io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [5:0]    io_read_2_cmd_payload,
  output wire [0:0]    io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [5:0]    io_read_3_cmd_payload,
  output wire [0:0]    io_read_3_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [0:0]    _zz_ram_0_port1;
  wire       [0:0]    _zz_ram_0_port2;
  wire       [0:0]    _zz_ram_0_port3;
  wire       [0:0]    _zz_ram_0_port4;
  wire       [0:0]    _zz_ram_0_port5;
  wire       [0:0]    _zz_ram_0_port6;
  wire       [0:0]    _zz_ram_0_port7;
  wire       [0:0]    _zz_ram_0_port8;
  wire       [0:0]    _zz_ram_0_port9;
  wire       [0:0]    _zz_ram_0_port10;
  wire       [0:0]    _zz_ram_0_port11;
  wire       [0:0]    _zz_ram_1_port0;
  wire       [0:0]    _zz_ram_1_port2;
  wire       [0:0]    _zz_ram_1_port3;
  wire       [0:0]    _zz_ram_1_port4;
  wire       [0:0]    _zz_ram_1_port5;
  wire       [0:0]    _zz_ram_1_port6;
  wire       [0:0]    _zz_ram_1_port7;
  wire       [0:0]    _zz_ram_1_port8;
  wire       [0:0]    _zz_ram_1_port9;
  wire       [0:0]    _zz_ram_1_port10;
  wire       [0:0]    _zz_ram_1_port11;
  wire       [0:0]    _zz_ram_2_port0;
  wire       [0:0]    _zz_ram_2_port1;
  wire       [0:0]    _zz_ram_2_port3;
  wire       [0:0]    _zz_ram_2_port4;
  wire       [0:0]    _zz_ram_2_port5;
  wire       [0:0]    _zz_ram_2_port6;
  wire       [0:0]    _zz_ram_2_port7;
  wire       [0:0]    _zz_ram_2_port8;
  wire       [0:0]    _zz_ram_2_port9;
  wire       [0:0]    _zz_ram_2_port10;
  wire       [0:0]    _zz_ram_2_port11;
  wire       [0:0]    _zz_ram_3_port0;
  wire       [0:0]    _zz_ram_3_port1;
  wire       [0:0]    _zz_ram_3_port2;
  wire       [0:0]    _zz_ram_3_port4;
  wire       [0:0]    _zz_ram_3_port5;
  wire       [0:0]    _zz_ram_3_port6;
  wire       [0:0]    _zz_ram_3_port7;
  wire       [0:0]    _zz_ram_3_port8;
  wire       [0:0]    _zz_ram_3_port9;
  wire       [0:0]    _zz_ram_3_port10;
  wire       [0:0]    _zz_ram_3_port11;
  wire       [0:0]    _zz_ram_4_port0;
  wire       [0:0]    _zz_ram_4_port1;
  wire       [0:0]    _zz_ram_4_port2;
  wire       [0:0]    _zz_ram_4_port3;
  wire       [0:0]    _zz_ram_4_port5;
  wire       [0:0]    _zz_ram_4_port6;
  wire       [0:0]    _zz_ram_4_port7;
  wire       [0:0]    _zz_ram_4_port8;
  wire       [0:0]    _zz_ram_4_port9;
  wire       [0:0]    _zz_ram_4_port10;
  wire       [0:0]    _zz_ram_4_port11;
  wire       [0:0]    _zz_ram_5_port0;
  wire       [0:0]    _zz_ram_5_port1;
  wire       [0:0]    _zz_ram_5_port2;
  wire       [0:0]    _zz_ram_5_port3;
  wire       [0:0]    _zz_ram_5_port4;
  wire       [0:0]    _zz_ram_5_port6;
  wire       [0:0]    _zz_ram_5_port7;
  wire       [0:0]    _zz_ram_5_port8;
  wire       [0:0]    _zz_ram_5_port9;
  wire       [0:0]    _zz_ram_5_port10;
  wire       [0:0]    _zz_ram_5_port11;
  wire       [0:0]    _zz_ram_6_port0;
  wire       [0:0]    _zz_ram_6_port1;
  wire       [0:0]    _zz_ram_6_port2;
  wire       [0:0]    _zz_ram_6_port3;
  wire       [0:0]    _zz_ram_6_port4;
  wire       [0:0]    _zz_ram_6_port5;
  wire       [0:0]    _zz_ram_6_port7;
  wire       [0:0]    _zz_ram_6_port8;
  wire       [0:0]    _zz_ram_6_port9;
  wire       [0:0]    _zz_ram_6_port10;
  wire       [0:0]    _zz_ram_6_port11;
  wire       [0:0]    _zz_ram_7_port0;
  wire       [0:0]    _zz_ram_7_port1;
  wire       [0:0]    _zz_ram_7_port2;
  wire       [0:0]    _zz_ram_7_port3;
  wire       [0:0]    _zz_ram_7_port4;
  wire       [0:0]    _zz_ram_7_port5;
  wire       [0:0]    _zz_ram_7_port6;
  wire       [0:0]    _zz_ram_7_port8;
  wire       [0:0]    _zz_ram_7_port9;
  wire       [0:0]    _zz_ram_7_port10;
  wire       [0:0]    _zz_ram_7_port11;
  wire       [0:0]    writes_0_values_0;
  wire       [0:0]    writes_0_values_1;
  wire       [0:0]    writes_0_values_2;
  wire       [0:0]    writes_0_values_3;
  wire       [0:0]    writes_0_values_4;
  wire       [0:0]    writes_0_values_5;
  wire       [0:0]    writes_0_values_6;
  wire       [0:0]    writes_0_xored;
  wire       [0:0]    writes_1_values_0;
  wire       [0:0]    writes_1_values_1;
  wire       [0:0]    writes_1_values_2;
  wire       [0:0]    writes_1_values_3;
  wire       [0:0]    writes_1_values_4;
  wire       [0:0]    writes_1_values_5;
  wire       [0:0]    writes_1_values_6;
  wire       [0:0]    writes_1_xored;
  wire       [0:0]    writes_2_values_0;
  wire       [0:0]    writes_2_values_1;
  wire       [0:0]    writes_2_values_2;
  wire       [0:0]    writes_2_values_3;
  wire       [0:0]    writes_2_values_4;
  wire       [0:0]    writes_2_values_5;
  wire       [0:0]    writes_2_values_6;
  wire       [0:0]    writes_2_xored;
  wire       [0:0]    writes_3_values_0;
  wire       [0:0]    writes_3_values_1;
  wire       [0:0]    writes_3_values_2;
  wire       [0:0]    writes_3_values_3;
  wire       [0:0]    writes_3_values_4;
  wire       [0:0]    writes_3_values_5;
  wire       [0:0]    writes_3_values_6;
  wire       [0:0]    writes_3_xored;
  wire       [0:0]    writes_4_values_0;
  wire       [0:0]    writes_4_values_1;
  wire       [0:0]    writes_4_values_2;
  wire       [0:0]    writes_4_values_3;
  wire       [0:0]    writes_4_values_4;
  wire       [0:0]    writes_4_values_5;
  wire       [0:0]    writes_4_values_6;
  wire       [0:0]    writes_4_xored;
  wire       [0:0]    writes_5_values_0;
  wire       [0:0]    writes_5_values_1;
  wire       [0:0]    writes_5_values_2;
  wire       [0:0]    writes_5_values_3;
  wire       [0:0]    writes_5_values_4;
  wire       [0:0]    writes_5_values_5;
  wire       [0:0]    writes_5_values_6;
  wire       [0:0]    writes_5_xored;
  wire       [0:0]    writes_6_values_0;
  wire       [0:0]    writes_6_values_1;
  wire       [0:0]    writes_6_values_2;
  wire       [0:0]    writes_6_values_3;
  wire       [0:0]    writes_6_values_4;
  wire       [0:0]    writes_6_values_5;
  wire       [0:0]    writes_6_values_6;
  wire       [0:0]    writes_6_xored;
  wire       [0:0]    writes_7_values_0;
  wire       [0:0]    writes_7_values_1;
  wire       [0:0]    writes_7_values_2;
  wire       [0:0]    writes_7_values_3;
  wire       [0:0]    writes_7_values_4;
  wire       [0:0]    writes_7_values_5;
  wire       [0:0]    writes_7_values_6;
  wire       [0:0]    writes_7_xored;
  wire       [0:0]    reads_0_values_0;
  wire       [0:0]    reads_0_values_1;
  wire       [0:0]    reads_0_values_2;
  wire       [0:0]    reads_0_values_3;
  wire       [0:0]    reads_0_values_4;
  wire       [0:0]    reads_0_values_5;
  wire       [0:0]    reads_0_values_6;
  wire       [0:0]    reads_0_values_7;
  wire       [0:0]    reads_0_xored;
  wire       [0:0]    reads_1_values_0;
  wire       [0:0]    reads_1_values_1;
  wire       [0:0]    reads_1_values_2;
  wire       [0:0]    reads_1_values_3;
  wire       [0:0]    reads_1_values_4;
  wire       [0:0]    reads_1_values_5;
  wire       [0:0]    reads_1_values_6;
  wire       [0:0]    reads_1_values_7;
  wire       [0:0]    reads_1_xored;
  wire       [0:0]    reads_2_values_0;
  wire       [0:0]    reads_2_values_1;
  wire       [0:0]    reads_2_values_2;
  wire       [0:0]    reads_2_values_3;
  wire       [0:0]    reads_2_values_4;
  wire       [0:0]    reads_2_values_5;
  wire       [0:0]    reads_2_values_6;
  wire       [0:0]    reads_2_values_7;
  wire       [0:0]    reads_2_xored;
  wire       [0:0]    reads_3_values_0;
  wire       [0:0]    reads_3_values_1;
  wire       [0:0]    reads_3_values_2;
  wire       [0:0]    reads_3_values_3;
  wire       [0:0]    reads_3_values_4;
  wire       [0:0]    reads_3_values_5;
  wire       [0:0]    reads_3_values_6;
  wire       [0:0]    reads_3_values_7;
  wire       [0:0]    reads_3_xored;
  (* ram_style = "distributed" *) reg [0:0] ram_0 [0:63];
  (* ram_style = "distributed" *) reg [0:0] ram_1 [0:63];
  (* ram_style = "distributed" *) reg [0:0] ram_2 [0:63];
  (* ram_style = "distributed" *) reg [0:0] ram_3 [0:63];
  (* ram_style = "distributed" *) reg [0:0] ram_4 [0:63];
  (* ram_style = "distributed" *) reg [0:0] ram_5 [0:63];
  (* ram_style = "distributed" *) reg [0:0] ram_6 [0:63];
  (* ram_style = "distributed" *) reg [0:0] ram_7 [0:63];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_writes_2_payload_address];
  assign _zz_ram_0_port3 = ram_0[io_writes_3_payload_address];
  assign _zz_ram_0_port4 = ram_0[io_writes_4_payload_address];
  assign _zz_ram_0_port5 = ram_0[io_writes_5_payload_address];
  assign _zz_ram_0_port6 = ram_0[io_writes_6_payload_address];
  assign _zz_ram_0_port7 = ram_0[io_writes_7_payload_address];
  assign _zz_ram_0_port8 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_0_port9 = ram_0[io_read_1_cmd_payload];
  assign _zz_ram_0_port10 = ram_0[io_read_2_cmd_payload];
  assign _zz_ram_0_port11 = ram_0[io_read_3_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_writes_2_payload_address];
  assign _zz_ram_1_port3 = ram_1[io_writes_3_payload_address];
  assign _zz_ram_1_port4 = ram_1[io_writes_4_payload_address];
  assign _zz_ram_1_port5 = ram_1[io_writes_5_payload_address];
  assign _zz_ram_1_port6 = ram_1[io_writes_6_payload_address];
  assign _zz_ram_1_port7 = ram_1[io_writes_7_payload_address];
  assign _zz_ram_1_port8 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_1_port9 = ram_1[io_read_1_cmd_payload];
  assign _zz_ram_1_port10 = ram_1[io_read_2_cmd_payload];
  assign _zz_ram_1_port11 = ram_1[io_read_3_cmd_payload];
  assign _zz_ram_2_port0 = ram_2[io_writes_0_payload_address];
  assign _zz_ram_2_port1 = ram_2[io_writes_1_payload_address];
  always @(posedge clk) begin
    if(io_writes_2_valid) begin
      ram_2[io_writes_2_payload_address] <= writes_2_xored;
    end
  end

  assign _zz_ram_2_port3 = ram_2[io_writes_3_payload_address];
  assign _zz_ram_2_port4 = ram_2[io_writes_4_payload_address];
  assign _zz_ram_2_port5 = ram_2[io_writes_5_payload_address];
  assign _zz_ram_2_port6 = ram_2[io_writes_6_payload_address];
  assign _zz_ram_2_port7 = ram_2[io_writes_7_payload_address];
  assign _zz_ram_2_port8 = ram_2[io_read_0_cmd_payload];
  assign _zz_ram_2_port9 = ram_2[io_read_1_cmd_payload];
  assign _zz_ram_2_port10 = ram_2[io_read_2_cmd_payload];
  assign _zz_ram_2_port11 = ram_2[io_read_3_cmd_payload];
  assign _zz_ram_3_port0 = ram_3[io_writes_0_payload_address];
  assign _zz_ram_3_port1 = ram_3[io_writes_1_payload_address];
  assign _zz_ram_3_port2 = ram_3[io_writes_2_payload_address];
  always @(posedge clk) begin
    if(io_writes_3_valid) begin
      ram_3[io_writes_3_payload_address] <= writes_3_xored;
    end
  end

  assign _zz_ram_3_port4 = ram_3[io_writes_4_payload_address];
  assign _zz_ram_3_port5 = ram_3[io_writes_5_payload_address];
  assign _zz_ram_3_port6 = ram_3[io_writes_6_payload_address];
  assign _zz_ram_3_port7 = ram_3[io_writes_7_payload_address];
  assign _zz_ram_3_port8 = ram_3[io_read_0_cmd_payload];
  assign _zz_ram_3_port9 = ram_3[io_read_1_cmd_payload];
  assign _zz_ram_3_port10 = ram_3[io_read_2_cmd_payload];
  assign _zz_ram_3_port11 = ram_3[io_read_3_cmd_payload];
  assign _zz_ram_4_port0 = ram_4[io_writes_0_payload_address];
  assign _zz_ram_4_port1 = ram_4[io_writes_1_payload_address];
  assign _zz_ram_4_port2 = ram_4[io_writes_2_payload_address];
  assign _zz_ram_4_port3 = ram_4[io_writes_3_payload_address];
  always @(posedge clk) begin
    if(io_writes_4_valid) begin
      ram_4[io_writes_4_payload_address] <= writes_4_xored;
    end
  end

  assign _zz_ram_4_port5 = ram_4[io_writes_5_payload_address];
  assign _zz_ram_4_port6 = ram_4[io_writes_6_payload_address];
  assign _zz_ram_4_port7 = ram_4[io_writes_7_payload_address];
  assign _zz_ram_4_port8 = ram_4[io_read_0_cmd_payload];
  assign _zz_ram_4_port9 = ram_4[io_read_1_cmd_payload];
  assign _zz_ram_4_port10 = ram_4[io_read_2_cmd_payload];
  assign _zz_ram_4_port11 = ram_4[io_read_3_cmd_payload];
  assign _zz_ram_5_port0 = ram_5[io_writes_0_payload_address];
  assign _zz_ram_5_port1 = ram_5[io_writes_1_payload_address];
  assign _zz_ram_5_port2 = ram_5[io_writes_2_payload_address];
  assign _zz_ram_5_port3 = ram_5[io_writes_3_payload_address];
  assign _zz_ram_5_port4 = ram_5[io_writes_4_payload_address];
  always @(posedge clk) begin
    if(io_writes_5_valid) begin
      ram_5[io_writes_5_payload_address] <= writes_5_xored;
    end
  end

  assign _zz_ram_5_port6 = ram_5[io_writes_6_payload_address];
  assign _zz_ram_5_port7 = ram_5[io_writes_7_payload_address];
  assign _zz_ram_5_port8 = ram_5[io_read_0_cmd_payload];
  assign _zz_ram_5_port9 = ram_5[io_read_1_cmd_payload];
  assign _zz_ram_5_port10 = ram_5[io_read_2_cmd_payload];
  assign _zz_ram_5_port11 = ram_5[io_read_3_cmd_payload];
  assign _zz_ram_6_port0 = ram_6[io_writes_0_payload_address];
  assign _zz_ram_6_port1 = ram_6[io_writes_1_payload_address];
  assign _zz_ram_6_port2 = ram_6[io_writes_2_payload_address];
  assign _zz_ram_6_port3 = ram_6[io_writes_3_payload_address];
  assign _zz_ram_6_port4 = ram_6[io_writes_4_payload_address];
  assign _zz_ram_6_port5 = ram_6[io_writes_5_payload_address];
  always @(posedge clk) begin
    if(io_writes_6_valid) begin
      ram_6[io_writes_6_payload_address] <= writes_6_xored;
    end
  end

  assign _zz_ram_6_port7 = ram_6[io_writes_7_payload_address];
  assign _zz_ram_6_port8 = ram_6[io_read_0_cmd_payload];
  assign _zz_ram_6_port9 = ram_6[io_read_1_cmd_payload];
  assign _zz_ram_6_port10 = ram_6[io_read_2_cmd_payload];
  assign _zz_ram_6_port11 = ram_6[io_read_3_cmd_payload];
  assign _zz_ram_7_port0 = ram_7[io_writes_0_payload_address];
  assign _zz_ram_7_port1 = ram_7[io_writes_1_payload_address];
  assign _zz_ram_7_port2 = ram_7[io_writes_2_payload_address];
  assign _zz_ram_7_port3 = ram_7[io_writes_3_payload_address];
  assign _zz_ram_7_port4 = ram_7[io_writes_4_payload_address];
  assign _zz_ram_7_port5 = ram_7[io_writes_5_payload_address];
  assign _zz_ram_7_port6 = ram_7[io_writes_6_payload_address];
  always @(posedge clk) begin
    if(io_writes_7_valid) begin
      ram_7[io_writes_7_payload_address] <= writes_7_xored;
    end
  end

  assign _zz_ram_7_port8 = ram_7[io_read_0_cmd_payload];
  assign _zz_ram_7_port9 = ram_7[io_read_1_cmd_payload];
  assign _zz_ram_7_port10 = ram_7[io_read_2_cmd_payload];
  assign _zz_ram_7_port11 = ram_7[io_read_3_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_values_1 = _zz_ram_2_port0;
  assign writes_0_values_2 = _zz_ram_3_port0;
  assign writes_0_values_3 = _zz_ram_4_port0;
  assign writes_0_values_4 = _zz_ram_5_port0;
  assign writes_0_values_5 = _zz_ram_6_port0;
  assign writes_0_values_6 = _zz_ram_7_port0;
  assign writes_0_xored = (((io_writes_0_payload_data ^ writes_0_values_0) ^ (writes_0_values_1 ^ writes_0_values_2)) ^ ((writes_0_values_3 ^ writes_0_values_4) ^ (writes_0_values_5 ^ writes_0_values_6)));
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_values_1 = _zz_ram_2_port1;
  assign writes_1_values_2 = _zz_ram_3_port1;
  assign writes_1_values_3 = _zz_ram_4_port1;
  assign writes_1_values_4 = _zz_ram_5_port1;
  assign writes_1_values_5 = _zz_ram_6_port1;
  assign writes_1_values_6 = _zz_ram_7_port1;
  assign writes_1_xored = (((io_writes_1_payload_data ^ writes_1_values_0) ^ (writes_1_values_1 ^ writes_1_values_2)) ^ ((writes_1_values_3 ^ writes_1_values_4) ^ (writes_1_values_5 ^ writes_1_values_6)));
  assign writes_2_values_0 = _zz_ram_0_port2;
  assign writes_2_values_1 = _zz_ram_1_port2;
  assign writes_2_values_2 = _zz_ram_3_port2;
  assign writes_2_values_3 = _zz_ram_4_port2;
  assign writes_2_values_4 = _zz_ram_5_port2;
  assign writes_2_values_5 = _zz_ram_6_port2;
  assign writes_2_values_6 = _zz_ram_7_port2;
  assign writes_2_xored = (((io_writes_2_payload_data ^ writes_2_values_0) ^ (writes_2_values_1 ^ writes_2_values_2)) ^ ((writes_2_values_3 ^ writes_2_values_4) ^ (writes_2_values_5 ^ writes_2_values_6)));
  assign writes_3_values_0 = _zz_ram_0_port3;
  assign writes_3_values_1 = _zz_ram_1_port3;
  assign writes_3_values_2 = _zz_ram_2_port3;
  assign writes_3_values_3 = _zz_ram_4_port3;
  assign writes_3_values_4 = _zz_ram_5_port3;
  assign writes_3_values_5 = _zz_ram_6_port3;
  assign writes_3_values_6 = _zz_ram_7_port3;
  assign writes_3_xored = (((io_writes_3_payload_data ^ writes_3_values_0) ^ (writes_3_values_1 ^ writes_3_values_2)) ^ ((writes_3_values_3 ^ writes_3_values_4) ^ (writes_3_values_5 ^ writes_3_values_6)));
  assign writes_4_values_0 = _zz_ram_0_port4;
  assign writes_4_values_1 = _zz_ram_1_port4;
  assign writes_4_values_2 = _zz_ram_2_port4;
  assign writes_4_values_3 = _zz_ram_3_port4;
  assign writes_4_values_4 = _zz_ram_5_port4;
  assign writes_4_values_5 = _zz_ram_6_port4;
  assign writes_4_values_6 = _zz_ram_7_port4;
  assign writes_4_xored = (((io_writes_4_payload_data ^ writes_4_values_0) ^ (writes_4_values_1 ^ writes_4_values_2)) ^ ((writes_4_values_3 ^ writes_4_values_4) ^ (writes_4_values_5 ^ writes_4_values_6)));
  assign writes_5_values_0 = _zz_ram_0_port5;
  assign writes_5_values_1 = _zz_ram_1_port5;
  assign writes_5_values_2 = _zz_ram_2_port5;
  assign writes_5_values_3 = _zz_ram_3_port5;
  assign writes_5_values_4 = _zz_ram_4_port5;
  assign writes_5_values_5 = _zz_ram_6_port5;
  assign writes_5_values_6 = _zz_ram_7_port5;
  assign writes_5_xored = (((io_writes_5_payload_data ^ writes_5_values_0) ^ (writes_5_values_1 ^ writes_5_values_2)) ^ ((writes_5_values_3 ^ writes_5_values_4) ^ (writes_5_values_5 ^ writes_5_values_6)));
  assign writes_6_values_0 = _zz_ram_0_port6;
  assign writes_6_values_1 = _zz_ram_1_port6;
  assign writes_6_values_2 = _zz_ram_2_port6;
  assign writes_6_values_3 = _zz_ram_3_port6;
  assign writes_6_values_4 = _zz_ram_4_port6;
  assign writes_6_values_5 = _zz_ram_5_port6;
  assign writes_6_values_6 = _zz_ram_7_port6;
  assign writes_6_xored = (((io_writes_6_payload_data ^ writes_6_values_0) ^ (writes_6_values_1 ^ writes_6_values_2)) ^ ((writes_6_values_3 ^ writes_6_values_4) ^ (writes_6_values_5 ^ writes_6_values_6)));
  assign writes_7_values_0 = _zz_ram_0_port7;
  assign writes_7_values_1 = _zz_ram_1_port7;
  assign writes_7_values_2 = _zz_ram_2_port7;
  assign writes_7_values_3 = _zz_ram_3_port7;
  assign writes_7_values_4 = _zz_ram_4_port7;
  assign writes_7_values_5 = _zz_ram_5_port7;
  assign writes_7_values_6 = _zz_ram_6_port7;
  assign writes_7_xored = (((io_writes_7_payload_data ^ writes_7_values_0) ^ (writes_7_values_1 ^ writes_7_values_2)) ^ ((writes_7_values_3 ^ writes_7_values_4) ^ (writes_7_values_5 ^ writes_7_values_6)));
  assign reads_0_values_0 = _zz_ram_0_port8;
  assign reads_0_values_1 = _zz_ram_1_port8;
  assign reads_0_values_2 = _zz_ram_2_port8;
  assign reads_0_values_3 = _zz_ram_3_port8;
  assign reads_0_values_4 = _zz_ram_4_port8;
  assign reads_0_values_5 = _zz_ram_5_port8;
  assign reads_0_values_6 = _zz_ram_6_port8;
  assign reads_0_values_7 = _zz_ram_7_port8;
  assign reads_0_xored = (((reads_0_values_0 ^ reads_0_values_1) ^ (reads_0_values_2 ^ reads_0_values_3)) ^ ((reads_0_values_4 ^ reads_0_values_5) ^ (reads_0_values_6 ^ reads_0_values_7)));
  assign io_read_0_rsp = reads_0_xored;
  assign reads_1_values_0 = _zz_ram_0_port9;
  assign reads_1_values_1 = _zz_ram_1_port9;
  assign reads_1_values_2 = _zz_ram_2_port9;
  assign reads_1_values_3 = _zz_ram_3_port9;
  assign reads_1_values_4 = _zz_ram_4_port9;
  assign reads_1_values_5 = _zz_ram_5_port9;
  assign reads_1_values_6 = _zz_ram_6_port9;
  assign reads_1_values_7 = _zz_ram_7_port9;
  assign reads_1_xored = (((reads_1_values_0 ^ reads_1_values_1) ^ (reads_1_values_2 ^ reads_1_values_3)) ^ ((reads_1_values_4 ^ reads_1_values_5) ^ (reads_1_values_6 ^ reads_1_values_7)));
  assign io_read_1_rsp = reads_1_xored;
  assign reads_2_values_0 = _zz_ram_0_port10;
  assign reads_2_values_1 = _zz_ram_1_port10;
  assign reads_2_values_2 = _zz_ram_2_port10;
  assign reads_2_values_3 = _zz_ram_3_port10;
  assign reads_2_values_4 = _zz_ram_4_port10;
  assign reads_2_values_5 = _zz_ram_5_port10;
  assign reads_2_values_6 = _zz_ram_6_port10;
  assign reads_2_values_7 = _zz_ram_7_port10;
  assign reads_2_xored = (((reads_2_values_0 ^ reads_2_values_1) ^ (reads_2_values_2 ^ reads_2_values_3)) ^ ((reads_2_values_4 ^ reads_2_values_5) ^ (reads_2_values_6 ^ reads_2_values_7)));
  assign io_read_2_rsp = reads_2_xored;
  assign reads_3_values_0 = _zz_ram_0_port11;
  assign reads_3_values_1 = _zz_ram_1_port11;
  assign reads_3_values_2 = _zz_ram_2_port11;
  assign reads_3_values_3 = _zz_ram_3_port11;
  assign reads_3_values_4 = _zz_ram_4_port11;
  assign reads_3_values_5 = _zz_ram_5_port11;
  assign reads_3_values_6 = _zz_ram_6_port11;
  assign reads_3_values_7 = _zz_ram_7_port11;
  assign reads_3_xored = (((reads_3_values_0 ^ reads_3_values_1) ^ (reads_3_values_2 ^ reads_3_values_3)) ^ ((reads_3_values_4 ^ reads_3_values_5) ^ (reads_3_values_6 ^ reads_3_values_7)));
  assign io_read_3_rsp = reads_3_xored;

endmodule

module RamAsyncMwXor_11 (
  input  wire          io_writes_0_valid,
  input  wire [5:0]    io_writes_0_payload_address,
  input  wire [5:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [5:0]    io_writes_1_payload_address,
  input  wire [5:0]    io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [5:0]    io_read_0_cmd_payload,
  output wire [5:0]    io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [5:0]    io_read_1_cmd_payload,
  output wire [5:0]    io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [5:0]    io_read_2_cmd_payload,
  output wire [5:0]    io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [5:0]    io_read_3_cmd_payload,
  output wire [5:0]    io_read_3_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [5:0]    _zz_ram_0_port1;
  wire       [5:0]    _zz_ram_0_port2;
  wire       [5:0]    _zz_ram_0_port3;
  wire       [5:0]    _zz_ram_0_port4;
  wire       [5:0]    _zz_ram_0_port5;
  wire       [5:0]    _zz_ram_1_port0;
  wire       [5:0]    _zz_ram_1_port2;
  wire       [5:0]    _zz_ram_1_port3;
  wire       [5:0]    _zz_ram_1_port4;
  wire       [5:0]    _zz_ram_1_port5;
  wire       [5:0]    writes_0_values_0;
  wire       [5:0]    writes_0_xored;
  wire       [5:0]    writes_1_values_0;
  wire       [5:0]    writes_1_xored;
  wire       [5:0]    reads_0_values_0;
  wire       [5:0]    reads_0_values_1;
  wire       [5:0]    reads_0_xored;
  wire       [5:0]    reads_1_values_0;
  wire       [5:0]    reads_1_values_1;
  wire       [5:0]    reads_1_xored;
  wire       [5:0]    reads_2_values_0;
  wire       [5:0]    reads_2_values_1;
  wire       [5:0]    reads_2_xored;
  wire       [5:0]    reads_3_values_0;
  wire       [5:0]    reads_3_values_1;
  wire       [5:0]    reads_3_xored;
  (* ram_style = "distributed" *) reg [5:0] ram_0 [0:63];
  (* ram_style = "distributed" *) reg [5:0] ram_1 [0:63];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_0_port3 = ram_0[io_read_1_cmd_payload];
  assign _zz_ram_0_port4 = ram_0[io_read_2_cmd_payload];
  assign _zz_ram_0_port5 = ram_0[io_read_3_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_1_port3 = ram_1[io_read_1_cmd_payload];
  assign _zz_ram_1_port4 = ram_1[io_read_2_cmd_payload];
  assign _zz_ram_1_port5 = ram_1[io_read_3_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_xored = (io_writes_0_payload_data ^ writes_0_values_0);
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_xored = (io_writes_1_payload_data ^ writes_1_values_0);
  assign reads_0_values_0 = _zz_ram_0_port2;
  assign reads_0_values_1 = _zz_ram_1_port2;
  assign reads_0_xored = (reads_0_values_0 ^ reads_0_values_1);
  assign io_read_0_rsp = reads_0_xored;
  assign reads_1_values_0 = _zz_ram_0_port3;
  assign reads_1_values_1 = _zz_ram_1_port3;
  assign reads_1_xored = (reads_1_values_0 ^ reads_1_values_1);
  assign io_read_1_rsp = reads_1_xored;
  assign reads_2_values_0 = _zz_ram_0_port4;
  assign reads_2_values_1 = _zz_ram_1_port4;
  assign reads_2_xored = (reads_2_values_0 ^ reads_2_values_1);
  assign io_read_2_rsp = reads_2_xored;
  assign reads_3_values_0 = _zz_ram_0_port5;
  assign reads_3_values_1 = _zz_ram_1_port5;
  assign reads_3_xored = (reads_3_values_0 ^ reads_3_values_1);
  assign io_read_3_rsp = reads_3_xored;

endmodule

module RamAsyncMwMux_3 (
  input  wire          io_writes_0_valid,
  input  wire [5:0]    io_writes_0_payload_address,
  input  wire [31:0]   io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [5:0]    io_writes_1_payload_address,
  input  wire [31:0]   io_writes_1_payload_data,
  input  wire          io_writes_2_valid,
  input  wire [5:0]    io_writes_2_payload_address,
  input  wire [31:0]   io_writes_2_payload_data,
  input  wire          io_writes_3_valid,
  input  wire [5:0]    io_writes_3_payload_address,
  input  wire [31:0]   io_writes_3_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [5:0]    io_read_0_cmd_payload,
  output wire [31:0]   io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [5:0]    io_read_1_cmd_payload,
  output wire [31:0]   io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [5:0]    io_read_2_cmd_payload,
  output wire [31:0]   io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [5:0]    io_read_3_cmd_payload,
  output wire [31:0]   io_read_3_rsp,
  input  wire          io_read_4_cmd_valid,
  input  wire [5:0]    io_read_4_cmd_payload,
  output wire [31:0]   io_read_4_rsp,
  input  wire          io_read_5_cmd_valid,
  input  wire [5:0]    io_read_5_cmd_payload,
  output wire [31:0]   io_read_5_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [1:0]    location_io_writes_0_payload_data;
  wire       [1:0]    location_io_writes_1_payload_data;
  wire       [1:0]    location_io_writes_2_payload_data;
  wire       [1:0]    location_io_writes_3_payload_data;
  wire       [31:0]   _zz_ram_0_port1;
  wire       [31:0]   _zz_ram_0_port2;
  wire       [31:0]   _zz_ram_0_port3;
  wire       [31:0]   _zz_ram_0_port4;
  wire       [31:0]   _zz_ram_0_port5;
  wire       [31:0]   _zz_ram_0_port6;
  wire       [31:0]   _zz_ram_1_port1;
  wire       [31:0]   _zz_ram_1_port2;
  wire       [31:0]   _zz_ram_1_port3;
  wire       [31:0]   _zz_ram_1_port4;
  wire       [31:0]   _zz_ram_1_port5;
  wire       [31:0]   _zz_ram_1_port6;
  wire       [31:0]   _zz_ram_2_port1;
  wire       [31:0]   _zz_ram_2_port2;
  wire       [31:0]   _zz_ram_2_port3;
  wire       [31:0]   _zz_ram_2_port4;
  wire       [31:0]   _zz_ram_2_port5;
  wire       [31:0]   _zz_ram_2_port6;
  wire       [31:0]   _zz_ram_3_port1;
  wire       [31:0]   _zz_ram_3_port2;
  wire       [31:0]   _zz_ram_3_port3;
  wire       [31:0]   _zz_ram_3_port4;
  wire       [31:0]   _zz_ram_3_port5;
  wire       [31:0]   _zz_ram_3_port6;
  wire       [1:0]    location_io_read_0_rsp;
  wire       [1:0]    location_io_read_1_rsp;
  wire       [1:0]    location_io_read_2_rsp;
  wire       [1:0]    location_io_read_3_rsp;
  wire       [1:0]    location_io_read_4_rsp;
  wire       [1:0]    location_io_read_5_rsp;
  reg        [31:0]   _zz_io_read_0_rsp;
  reg        [31:0]   _zz_io_read_1_rsp;
  reg        [31:0]   _zz_io_read_2_rsp;
  reg        [31:0]   _zz_io_read_3_rsp;
  reg        [31:0]   _zz_io_read_4_rsp;
  reg        [31:0]   _zz_io_read_5_rsp;
  wire       [31:0]   reads_0_reads_0;
  wire       [31:0]   reads_0_reads_1;
  wire       [31:0]   reads_0_reads_2;
  wire       [31:0]   reads_0_reads_3;
  wire       [31:0]   reads_1_reads_0;
  wire       [31:0]   reads_1_reads_1;
  wire       [31:0]   reads_1_reads_2;
  wire       [31:0]   reads_1_reads_3;
  wire       [31:0]   reads_2_reads_0;
  wire       [31:0]   reads_2_reads_1;
  wire       [31:0]   reads_2_reads_2;
  wire       [31:0]   reads_2_reads_3;
  wire       [31:0]   reads_3_reads_0;
  wire       [31:0]   reads_3_reads_1;
  wire       [31:0]   reads_3_reads_2;
  wire       [31:0]   reads_3_reads_3;
  wire       [31:0]   reads_4_reads_0;
  wire       [31:0]   reads_4_reads_1;
  wire       [31:0]   reads_4_reads_2;
  wire       [31:0]   reads_4_reads_3;
  wire       [31:0]   reads_5_reads_0;
  wire       [31:0]   reads_5_reads_1;
  wire       [31:0]   reads_5_reads_2;
  wire       [31:0]   reads_5_reads_3;
  (* ram_style = "distributed" *) reg [31:0] ram_0 [0:63] /* verilator public */ ;
  (* ram_style = "distributed" *) reg [31:0] ram_1 [0:63] /* verilator public */ ;
  (* ram_style = "distributed" *) reg [31:0] ram_2 [0:63] /* verilator public */ ;
  (* ram_style = "distributed" *) reg [31:0] ram_3 [0:63] /* verilator public */ ;

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= io_writes_0_payload_data;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_0_port2 = ram_0[io_read_1_cmd_payload];
  assign _zz_ram_0_port3 = ram_0[io_read_2_cmd_payload];
  assign _zz_ram_0_port4 = ram_0[io_read_3_cmd_payload];
  assign _zz_ram_0_port5 = ram_0[io_read_4_cmd_payload];
  assign _zz_ram_0_port6 = ram_0[io_read_5_cmd_payload];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= io_writes_1_payload_data;
    end
  end

  assign _zz_ram_1_port1 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_1_port2 = ram_1[io_read_1_cmd_payload];
  assign _zz_ram_1_port3 = ram_1[io_read_2_cmd_payload];
  assign _zz_ram_1_port4 = ram_1[io_read_3_cmd_payload];
  assign _zz_ram_1_port5 = ram_1[io_read_4_cmd_payload];
  assign _zz_ram_1_port6 = ram_1[io_read_5_cmd_payload];
  always @(posedge clk) begin
    if(io_writes_2_valid) begin
      ram_2[io_writes_2_payload_address] <= io_writes_2_payload_data;
    end
  end

  assign _zz_ram_2_port1 = ram_2[io_read_0_cmd_payload];
  assign _zz_ram_2_port2 = ram_2[io_read_1_cmd_payload];
  assign _zz_ram_2_port3 = ram_2[io_read_2_cmd_payload];
  assign _zz_ram_2_port4 = ram_2[io_read_3_cmd_payload];
  assign _zz_ram_2_port5 = ram_2[io_read_4_cmd_payload];
  assign _zz_ram_2_port6 = ram_2[io_read_5_cmd_payload];
  always @(posedge clk) begin
    if(io_writes_3_valid) begin
      ram_3[io_writes_3_payload_address] <= io_writes_3_payload_data;
    end
  end

  assign _zz_ram_3_port1 = ram_3[io_read_0_cmd_payload];
  assign _zz_ram_3_port2 = ram_3[io_read_1_cmd_payload];
  assign _zz_ram_3_port3 = ram_3[io_read_2_cmd_payload];
  assign _zz_ram_3_port4 = ram_3[io_read_3_cmd_payload];
  assign _zz_ram_3_port5 = ram_3[io_read_4_cmd_payload];
  assign _zz_ram_3_port6 = ram_3[io_read_5_cmd_payload];
  RamAsyncMwXor_15 location (
    .io_writes_0_valid           (io_writes_0_valid                     ), //i
    .io_writes_0_payload_address (io_writes_0_payload_address[5:0]      ), //i
    .io_writes_0_payload_data    (location_io_writes_0_payload_data[1:0]), //i
    .io_writes_1_valid           (io_writes_1_valid                     ), //i
    .io_writes_1_payload_address (io_writes_1_payload_address[5:0]      ), //i
    .io_writes_1_payload_data    (location_io_writes_1_payload_data[1:0]), //i
    .io_writes_2_valid           (io_writes_2_valid                     ), //i
    .io_writes_2_payload_address (io_writes_2_payload_address[5:0]      ), //i
    .io_writes_2_payload_data    (location_io_writes_2_payload_data[1:0]), //i
    .io_writes_3_valid           (io_writes_3_valid                     ), //i
    .io_writes_3_payload_address (io_writes_3_payload_address[5:0]      ), //i
    .io_writes_3_payload_data    (location_io_writes_3_payload_data[1:0]), //i
    .io_read_0_cmd_valid         (io_read_0_cmd_valid                   ), //i
    .io_read_0_cmd_payload       (io_read_0_cmd_payload[5:0]            ), //i
    .io_read_0_rsp               (location_io_read_0_rsp[1:0]           ), //o
    .io_read_1_cmd_valid         (io_read_1_cmd_valid                   ), //i
    .io_read_1_cmd_payload       (io_read_1_cmd_payload[5:0]            ), //i
    .io_read_1_rsp               (location_io_read_1_rsp[1:0]           ), //o
    .io_read_2_cmd_valid         (io_read_2_cmd_valid                   ), //i
    .io_read_2_cmd_payload       (io_read_2_cmd_payload[5:0]            ), //i
    .io_read_2_rsp               (location_io_read_2_rsp[1:0]           ), //o
    .io_read_3_cmd_valid         (io_read_3_cmd_valid                   ), //i
    .io_read_3_cmd_payload       (io_read_3_cmd_payload[5:0]            ), //i
    .io_read_3_rsp               (location_io_read_3_rsp[1:0]           ), //o
    .io_read_4_cmd_valid         (io_read_4_cmd_valid                   ), //i
    .io_read_4_cmd_payload       (io_read_4_cmd_payload[5:0]            ), //i
    .io_read_4_rsp               (location_io_read_4_rsp[1:0]           ), //o
    .io_read_5_cmd_valid         (io_read_5_cmd_valid                   ), //i
    .io_read_5_cmd_payload       (io_read_5_cmd_payload[5:0]            ), //i
    .io_read_5_rsp               (location_io_read_5_rsp[1:0]           ), //o
    .clk                         (clk                                   ), //i
    .reset                       (reset                                 )  //i
  );
  always @(*) begin
    case(location_io_read_0_rsp)
      2'b00 : _zz_io_read_0_rsp = reads_0_reads_0;
      2'b01 : _zz_io_read_0_rsp = reads_0_reads_1;
      2'b10 : _zz_io_read_0_rsp = reads_0_reads_2;
      default : _zz_io_read_0_rsp = reads_0_reads_3;
    endcase
  end

  always @(*) begin
    case(location_io_read_1_rsp)
      2'b00 : _zz_io_read_1_rsp = reads_1_reads_0;
      2'b01 : _zz_io_read_1_rsp = reads_1_reads_1;
      2'b10 : _zz_io_read_1_rsp = reads_1_reads_2;
      default : _zz_io_read_1_rsp = reads_1_reads_3;
    endcase
  end

  always @(*) begin
    case(location_io_read_2_rsp)
      2'b00 : _zz_io_read_2_rsp = reads_2_reads_0;
      2'b01 : _zz_io_read_2_rsp = reads_2_reads_1;
      2'b10 : _zz_io_read_2_rsp = reads_2_reads_2;
      default : _zz_io_read_2_rsp = reads_2_reads_3;
    endcase
  end

  always @(*) begin
    case(location_io_read_3_rsp)
      2'b00 : _zz_io_read_3_rsp = reads_3_reads_0;
      2'b01 : _zz_io_read_3_rsp = reads_3_reads_1;
      2'b10 : _zz_io_read_3_rsp = reads_3_reads_2;
      default : _zz_io_read_3_rsp = reads_3_reads_3;
    endcase
  end

  always @(*) begin
    case(location_io_read_4_rsp)
      2'b00 : _zz_io_read_4_rsp = reads_4_reads_0;
      2'b01 : _zz_io_read_4_rsp = reads_4_reads_1;
      2'b10 : _zz_io_read_4_rsp = reads_4_reads_2;
      default : _zz_io_read_4_rsp = reads_4_reads_3;
    endcase
  end

  always @(*) begin
    case(location_io_read_5_rsp)
      2'b00 : _zz_io_read_5_rsp = reads_5_reads_0;
      2'b01 : _zz_io_read_5_rsp = reads_5_reads_1;
      2'b10 : _zz_io_read_5_rsp = reads_5_reads_2;
      default : _zz_io_read_5_rsp = reads_5_reads_3;
    endcase
  end

  assign location_io_writes_0_payload_data = 2'b00;
  assign location_io_writes_1_payload_data = 2'b01;
  assign location_io_writes_2_payload_data = 2'b10;
  assign location_io_writes_3_payload_data = 2'b11;
  assign reads_0_reads_0 = _zz_ram_0_port1;
  assign reads_0_reads_1 = _zz_ram_1_port1;
  assign reads_0_reads_2 = _zz_ram_2_port1;
  assign reads_0_reads_3 = _zz_ram_3_port1;
  assign io_read_0_rsp = _zz_io_read_0_rsp;
  assign reads_1_reads_0 = _zz_ram_0_port2;
  assign reads_1_reads_1 = _zz_ram_1_port2;
  assign reads_1_reads_2 = _zz_ram_2_port2;
  assign reads_1_reads_3 = _zz_ram_3_port2;
  assign io_read_1_rsp = _zz_io_read_1_rsp;
  assign reads_2_reads_0 = _zz_ram_0_port3;
  assign reads_2_reads_1 = _zz_ram_1_port3;
  assign reads_2_reads_2 = _zz_ram_2_port3;
  assign reads_2_reads_3 = _zz_ram_3_port3;
  assign io_read_2_rsp = _zz_io_read_2_rsp;
  assign reads_3_reads_0 = _zz_ram_0_port4;
  assign reads_3_reads_1 = _zz_ram_1_port4;
  assign reads_3_reads_2 = _zz_ram_2_port4;
  assign reads_3_reads_3 = _zz_ram_3_port4;
  assign io_read_3_rsp = _zz_io_read_3_rsp;
  assign reads_4_reads_0 = _zz_ram_0_port5;
  assign reads_4_reads_1 = _zz_ram_1_port5;
  assign reads_4_reads_2 = _zz_ram_2_port5;
  assign reads_4_reads_3 = _zz_ram_3_port5;
  assign io_read_4_rsp = _zz_io_read_4_rsp;
  assign reads_5_reads_0 = _zz_ram_0_port6;
  assign reads_5_reads_1 = _zz_ram_1_port6;
  assign reads_5_reads_2 = _zz_ram_2_port6;
  assign reads_5_reads_3 = _zz_ram_3_port6;
  assign io_read_5_rsp = _zz_io_read_5_rsp;

endmodule

module StreamFifo (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [5:0]    io_push_payload_robId,
  input  wire [1:0]    io_push_payload_mask,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [5:0]    io_pop_payload_robId,
  output wire [1:0]    io_pop_payload_mask,
  input  wire          io_flush,
  output wire [5:0]    io_occupancy,
  output wire [5:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  wire       [7:0]    _zz_logic_ram_port1;
  wire       [7:0]    _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [5:0]    logic_ptr_push;
  reg        [5:0]    logic_ptr_pop;
  wire       [5:0]    logic_ptr_occupancy;
  wire       [5:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1205;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [4:0]    logic_push_onRam_write_payload_address;
  wire       [5:0]    logic_push_onRam_write_payload_data_robId;
  wire       [1:0]    logic_push_onRam_write_payload_data_mask;
  wire                logic_pop_addressGen_valid;
  wire                logic_pop_addressGen_ready;
  wire       [4:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire       [5:0]    logic_pop_async_readed_robId;
  wire       [1:0]    logic_pop_async_readed_mask;
  wire       [7:0]    _zz_logic_pop_async_readed_robId;
  wire                logic_pop_addressGen_translated_valid;
  wire                logic_pop_addressGen_translated_ready;
  wire       [5:0]    logic_pop_addressGen_translated_payload_robId;
  wire       [1:0]    logic_pop_addressGen_translated_payload_mask;
  (* ram_style = "distributed" *) reg [7:0] logic_ram [0:31];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_mask,logic_push_onRam_write_payload_data_robId};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  assign _zz_logic_ram_port1 = logic_ram[logic_pop_addressGen_payload];
  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1205 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 6'h20) == 6'h00);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[4:0];
  assign logic_push_onRam_write_payload_data_robId = io_push_payload_robId;
  assign logic_push_onRam_write_payload_data_mask = io_push_payload_mask;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[4:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  assign _zz_logic_pop_async_readed_robId = _zz_logic_ram_port1;
  assign logic_pop_async_readed_robId = _zz_logic_pop_async_readed_robId[5 : 0];
  assign logic_pop_async_readed_mask = _zz_logic_pop_async_readed_robId[7 : 6];
  assign logic_pop_addressGen_translated_valid = logic_pop_addressGen_valid;
  assign logic_pop_addressGen_ready = logic_pop_addressGen_translated_ready;
  assign logic_pop_addressGen_translated_payload_robId = logic_pop_async_readed_robId;
  assign logic_pop_addressGen_translated_payload_mask = logic_pop_async_readed_mask;
  assign io_pop_valid = logic_pop_addressGen_translated_valid;
  assign logic_pop_addressGen_translated_ready = io_pop_ready;
  assign io_pop_payload_robId = logic_pop_addressGen_translated_payload_robId;
  assign io_pop_payload_mask = logic_pop_addressGen_translated_payload_mask;
  assign logic_ptr_popOnIo = logic_ptr_pop;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (6'h20 - logic_ptr_occupancy);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      logic_ptr_push <= 6'h00;
      logic_ptr_pop <= 6'h00;
      logic_ptr_wentUp <= 1'b0;
    end else begin
      if(when_Stream_l1205) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 6'h01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 6'h01);
      end
      if(io_flush) begin
        logic_ptr_push <= 6'h00;
        logic_ptr_pop <= 6'h00;
      end
    end
  end


endmodule

//RamAsyncMwXor_14 replaced by RamAsyncMwXor_13

module RamAsyncMwXor_13 (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_payload_address,
  input  wire [5:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [4:0]    io_writes_1_payload_address,
  input  wire [5:0]    io_writes_1_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [4:0]    io_read_0_cmd_payload,
  output wire [5:0]    io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [4:0]    io_read_1_cmd_payload,
  output wire [5:0]    io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [4:0]    io_read_2_cmd_payload,
  output wire [5:0]    io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [4:0]    io_read_3_cmd_payload,
  output wire [5:0]    io_read_3_rsp,
  input  wire          io_read_4_cmd_valid,
  input  wire [4:0]    io_read_4_cmd_payload,
  output wire [5:0]    io_read_4_rsp,
  input  wire          io_read_5_cmd_valid,
  input  wire [4:0]    io_read_5_cmd_payload,
  output wire [5:0]    io_read_5_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [5:0]    _zz_ram_0_port1;
  wire       [5:0]    _zz_ram_0_port2;
  wire       [5:0]    _zz_ram_0_port3;
  wire       [5:0]    _zz_ram_0_port4;
  wire       [5:0]    _zz_ram_0_port5;
  wire       [5:0]    _zz_ram_0_port6;
  wire       [5:0]    _zz_ram_0_port7;
  wire       [5:0]    _zz_ram_1_port0;
  wire       [5:0]    _zz_ram_1_port2;
  wire       [5:0]    _zz_ram_1_port3;
  wire       [5:0]    _zz_ram_1_port4;
  wire       [5:0]    _zz_ram_1_port5;
  wire       [5:0]    _zz_ram_1_port6;
  wire       [5:0]    _zz_ram_1_port7;
  wire       [5:0]    writes_0_values_0;
  wire       [5:0]    writes_0_xored;
  wire       [5:0]    writes_1_values_0;
  wire       [5:0]    writes_1_xored;
  wire       [5:0]    reads_0_values_0;
  wire       [5:0]    reads_0_values_1;
  wire       [5:0]    reads_0_xored;
  wire       [5:0]    reads_1_values_0;
  wire       [5:0]    reads_1_values_1;
  wire       [5:0]    reads_1_xored;
  wire       [5:0]    reads_2_values_0;
  wire       [5:0]    reads_2_values_1;
  wire       [5:0]    reads_2_xored;
  wire       [5:0]    reads_3_values_0;
  wire       [5:0]    reads_3_values_1;
  wire       [5:0]    reads_3_xored;
  wire       [5:0]    reads_4_values_0;
  wire       [5:0]    reads_4_values_1;
  wire       [5:0]    reads_4_xored;
  wire       [5:0]    reads_5_values_0;
  wire       [5:0]    reads_5_values_1;
  wire       [5:0]    reads_5_xored;
  (* ram_style = "distributed" *) reg [5:0] ram_0 [0:31];
  (* ram_style = "distributed" *) reg [5:0] ram_1 [0:31];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_0_port3 = ram_0[io_read_1_cmd_payload];
  assign _zz_ram_0_port4 = ram_0[io_read_2_cmd_payload];
  assign _zz_ram_0_port5 = ram_0[io_read_3_cmd_payload];
  assign _zz_ram_0_port6 = ram_0[io_read_4_cmd_payload];
  assign _zz_ram_0_port7 = ram_0[io_read_5_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_1_port3 = ram_1[io_read_1_cmd_payload];
  assign _zz_ram_1_port4 = ram_1[io_read_2_cmd_payload];
  assign _zz_ram_1_port5 = ram_1[io_read_3_cmd_payload];
  assign _zz_ram_1_port6 = ram_1[io_read_4_cmd_payload];
  assign _zz_ram_1_port7 = ram_1[io_read_5_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_xored = (io_writes_0_payload_data ^ writes_0_values_0);
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_xored = (io_writes_1_payload_data ^ writes_1_values_0);
  assign reads_0_values_0 = _zz_ram_0_port2;
  assign reads_0_values_1 = _zz_ram_1_port2;
  assign reads_0_xored = (reads_0_values_0 ^ reads_0_values_1);
  assign io_read_0_rsp = reads_0_xored;
  assign reads_1_values_0 = _zz_ram_0_port3;
  assign reads_1_values_1 = _zz_ram_1_port3;
  assign reads_1_xored = (reads_1_values_0 ^ reads_1_values_1);
  assign io_read_1_rsp = reads_1_xored;
  assign reads_2_values_0 = _zz_ram_0_port4;
  assign reads_2_values_1 = _zz_ram_1_port4;
  assign reads_2_xored = (reads_2_values_0 ^ reads_2_values_1);
  assign io_read_2_rsp = reads_2_xored;
  assign reads_3_values_0 = _zz_ram_0_port5;
  assign reads_3_values_1 = _zz_ram_1_port5;
  assign reads_3_xored = (reads_3_values_0 ^ reads_3_values_1);
  assign io_read_3_rsp = reads_3_xored;
  assign reads_4_values_0 = _zz_ram_0_port6;
  assign reads_4_values_1 = _zz_ram_1_port6;
  assign reads_4_xored = (reads_4_values_0 ^ reads_4_values_1);
  assign io_read_4_rsp = reads_4_xored;
  assign reads_5_values_0 = _zz_ram_0_port7;
  assign reads_5_values_1 = _zz_ram_1_port7;
  assign reads_5_xored = (reads_5_values_0 ^ reads_5_values_1);
  assign io_read_5_rsp = reads_5_xored;

endmodule

module RamAsyncMwXor_15 (
  input  wire          io_writes_0_valid,
  input  wire [5:0]    io_writes_0_payload_address,
  input  wire [1:0]    io_writes_0_payload_data,
  input  wire          io_writes_1_valid,
  input  wire [5:0]    io_writes_1_payload_address,
  input  wire [1:0]    io_writes_1_payload_data,
  input  wire          io_writes_2_valid,
  input  wire [5:0]    io_writes_2_payload_address,
  input  wire [1:0]    io_writes_2_payload_data,
  input  wire          io_writes_3_valid,
  input  wire [5:0]    io_writes_3_payload_address,
  input  wire [1:0]    io_writes_3_payload_data,
  input  wire          io_read_0_cmd_valid,
  input  wire [5:0]    io_read_0_cmd_payload,
  output wire [1:0]    io_read_0_rsp,
  input  wire          io_read_1_cmd_valid,
  input  wire [5:0]    io_read_1_cmd_payload,
  output wire [1:0]    io_read_1_rsp,
  input  wire          io_read_2_cmd_valid,
  input  wire [5:0]    io_read_2_cmd_payload,
  output wire [1:0]    io_read_2_rsp,
  input  wire          io_read_3_cmd_valid,
  input  wire [5:0]    io_read_3_cmd_payload,
  output wire [1:0]    io_read_3_rsp,
  input  wire          io_read_4_cmd_valid,
  input  wire [5:0]    io_read_4_cmd_payload,
  output wire [1:0]    io_read_4_rsp,
  input  wire          io_read_5_cmd_valid,
  input  wire [5:0]    io_read_5_cmd_payload,
  output wire [1:0]    io_read_5_rsp,
  input  wire          clk,
  input  wire          reset
);

  wire       [1:0]    _zz_ram_0_port1;
  wire       [1:0]    _zz_ram_0_port2;
  wire       [1:0]    _zz_ram_0_port3;
  wire       [1:0]    _zz_ram_0_port4;
  wire       [1:0]    _zz_ram_0_port5;
  wire       [1:0]    _zz_ram_0_port6;
  wire       [1:0]    _zz_ram_0_port7;
  wire       [1:0]    _zz_ram_0_port8;
  wire       [1:0]    _zz_ram_0_port9;
  wire       [1:0]    _zz_ram_1_port0;
  wire       [1:0]    _zz_ram_1_port2;
  wire       [1:0]    _zz_ram_1_port3;
  wire       [1:0]    _zz_ram_1_port4;
  wire       [1:0]    _zz_ram_1_port5;
  wire       [1:0]    _zz_ram_1_port6;
  wire       [1:0]    _zz_ram_1_port7;
  wire       [1:0]    _zz_ram_1_port8;
  wire       [1:0]    _zz_ram_1_port9;
  wire       [1:0]    _zz_ram_2_port0;
  wire       [1:0]    _zz_ram_2_port1;
  wire       [1:0]    _zz_ram_2_port3;
  wire       [1:0]    _zz_ram_2_port4;
  wire       [1:0]    _zz_ram_2_port5;
  wire       [1:0]    _zz_ram_2_port6;
  wire       [1:0]    _zz_ram_2_port7;
  wire       [1:0]    _zz_ram_2_port8;
  wire       [1:0]    _zz_ram_2_port9;
  wire       [1:0]    _zz_ram_3_port0;
  wire       [1:0]    _zz_ram_3_port1;
  wire       [1:0]    _zz_ram_3_port2;
  wire       [1:0]    _zz_ram_3_port4;
  wire       [1:0]    _zz_ram_3_port5;
  wire       [1:0]    _zz_ram_3_port6;
  wire       [1:0]    _zz_ram_3_port7;
  wire       [1:0]    _zz_ram_3_port8;
  wire       [1:0]    _zz_ram_3_port9;
  wire       [1:0]    writes_0_values_0;
  wire       [1:0]    writes_0_values_1;
  wire       [1:0]    writes_0_values_2;
  wire       [1:0]    writes_0_xored;
  wire       [1:0]    writes_1_values_0;
  wire       [1:0]    writes_1_values_1;
  wire       [1:0]    writes_1_values_2;
  wire       [1:0]    writes_1_xored;
  wire       [1:0]    writes_2_values_0;
  wire       [1:0]    writes_2_values_1;
  wire       [1:0]    writes_2_values_2;
  wire       [1:0]    writes_2_xored;
  wire       [1:0]    writes_3_values_0;
  wire       [1:0]    writes_3_values_1;
  wire       [1:0]    writes_3_values_2;
  wire       [1:0]    writes_3_xored;
  wire       [1:0]    reads_0_values_0;
  wire       [1:0]    reads_0_values_1;
  wire       [1:0]    reads_0_values_2;
  wire       [1:0]    reads_0_values_3;
  wire       [1:0]    reads_0_xored;
  wire       [1:0]    reads_1_values_0;
  wire       [1:0]    reads_1_values_1;
  wire       [1:0]    reads_1_values_2;
  wire       [1:0]    reads_1_values_3;
  wire       [1:0]    reads_1_xored;
  wire       [1:0]    reads_2_values_0;
  wire       [1:0]    reads_2_values_1;
  wire       [1:0]    reads_2_values_2;
  wire       [1:0]    reads_2_values_3;
  wire       [1:0]    reads_2_xored;
  wire       [1:0]    reads_3_values_0;
  wire       [1:0]    reads_3_values_1;
  wire       [1:0]    reads_3_values_2;
  wire       [1:0]    reads_3_values_3;
  wire       [1:0]    reads_3_xored;
  wire       [1:0]    reads_4_values_0;
  wire       [1:0]    reads_4_values_1;
  wire       [1:0]    reads_4_values_2;
  wire       [1:0]    reads_4_values_3;
  wire       [1:0]    reads_4_xored;
  wire       [1:0]    reads_5_values_0;
  wire       [1:0]    reads_5_values_1;
  wire       [1:0]    reads_5_values_2;
  wire       [1:0]    reads_5_values_3;
  wire       [1:0]    reads_5_xored;
  (* ram_style = "distributed" *) reg [1:0] ram_0 [0:63];
  (* ram_style = "distributed" *) reg [1:0] ram_1 [0:63];
  (* ram_style = "distributed" *) reg [1:0] ram_2 [0:63];
  (* ram_style = "distributed" *) reg [1:0] ram_3 [0:63];

  always @(posedge clk) begin
    if(io_writes_0_valid) begin
      ram_0[io_writes_0_payload_address] <= writes_0_xored;
    end
  end

  assign _zz_ram_0_port1 = ram_0[io_writes_1_payload_address];
  assign _zz_ram_0_port2 = ram_0[io_writes_2_payload_address];
  assign _zz_ram_0_port3 = ram_0[io_writes_3_payload_address];
  assign _zz_ram_0_port4 = ram_0[io_read_0_cmd_payload];
  assign _zz_ram_0_port5 = ram_0[io_read_1_cmd_payload];
  assign _zz_ram_0_port6 = ram_0[io_read_2_cmd_payload];
  assign _zz_ram_0_port7 = ram_0[io_read_3_cmd_payload];
  assign _zz_ram_0_port8 = ram_0[io_read_4_cmd_payload];
  assign _zz_ram_0_port9 = ram_0[io_read_5_cmd_payload];
  assign _zz_ram_1_port0 = ram_1[io_writes_0_payload_address];
  always @(posedge clk) begin
    if(io_writes_1_valid) begin
      ram_1[io_writes_1_payload_address] <= writes_1_xored;
    end
  end

  assign _zz_ram_1_port2 = ram_1[io_writes_2_payload_address];
  assign _zz_ram_1_port3 = ram_1[io_writes_3_payload_address];
  assign _zz_ram_1_port4 = ram_1[io_read_0_cmd_payload];
  assign _zz_ram_1_port5 = ram_1[io_read_1_cmd_payload];
  assign _zz_ram_1_port6 = ram_1[io_read_2_cmd_payload];
  assign _zz_ram_1_port7 = ram_1[io_read_3_cmd_payload];
  assign _zz_ram_1_port8 = ram_1[io_read_4_cmd_payload];
  assign _zz_ram_1_port9 = ram_1[io_read_5_cmd_payload];
  assign _zz_ram_2_port0 = ram_2[io_writes_0_payload_address];
  assign _zz_ram_2_port1 = ram_2[io_writes_1_payload_address];
  always @(posedge clk) begin
    if(io_writes_2_valid) begin
      ram_2[io_writes_2_payload_address] <= writes_2_xored;
    end
  end

  assign _zz_ram_2_port3 = ram_2[io_writes_3_payload_address];
  assign _zz_ram_2_port4 = ram_2[io_read_0_cmd_payload];
  assign _zz_ram_2_port5 = ram_2[io_read_1_cmd_payload];
  assign _zz_ram_2_port6 = ram_2[io_read_2_cmd_payload];
  assign _zz_ram_2_port7 = ram_2[io_read_3_cmd_payload];
  assign _zz_ram_2_port8 = ram_2[io_read_4_cmd_payload];
  assign _zz_ram_2_port9 = ram_2[io_read_5_cmd_payload];
  assign _zz_ram_3_port0 = ram_3[io_writes_0_payload_address];
  assign _zz_ram_3_port1 = ram_3[io_writes_1_payload_address];
  assign _zz_ram_3_port2 = ram_3[io_writes_2_payload_address];
  always @(posedge clk) begin
    if(io_writes_3_valid) begin
      ram_3[io_writes_3_payload_address] <= writes_3_xored;
    end
  end

  assign _zz_ram_3_port4 = ram_3[io_read_0_cmd_payload];
  assign _zz_ram_3_port5 = ram_3[io_read_1_cmd_payload];
  assign _zz_ram_3_port6 = ram_3[io_read_2_cmd_payload];
  assign _zz_ram_3_port7 = ram_3[io_read_3_cmd_payload];
  assign _zz_ram_3_port8 = ram_3[io_read_4_cmd_payload];
  assign _zz_ram_3_port9 = ram_3[io_read_5_cmd_payload];
  assign writes_0_values_0 = _zz_ram_1_port0;
  assign writes_0_values_1 = _zz_ram_2_port0;
  assign writes_0_values_2 = _zz_ram_3_port0;
  assign writes_0_xored = ((io_writes_0_payload_data ^ writes_0_values_0) ^ (writes_0_values_1 ^ writes_0_values_2));
  assign writes_1_values_0 = _zz_ram_0_port1;
  assign writes_1_values_1 = _zz_ram_2_port1;
  assign writes_1_values_2 = _zz_ram_3_port1;
  assign writes_1_xored = ((io_writes_1_payload_data ^ writes_1_values_0) ^ (writes_1_values_1 ^ writes_1_values_2));
  assign writes_2_values_0 = _zz_ram_0_port2;
  assign writes_2_values_1 = _zz_ram_1_port2;
  assign writes_2_values_2 = _zz_ram_3_port2;
  assign writes_2_xored = ((io_writes_2_payload_data ^ writes_2_values_0) ^ (writes_2_values_1 ^ writes_2_values_2));
  assign writes_3_values_0 = _zz_ram_0_port3;
  assign writes_3_values_1 = _zz_ram_1_port3;
  assign writes_3_values_2 = _zz_ram_2_port3;
  assign writes_3_xored = ((io_writes_3_payload_data ^ writes_3_values_0) ^ (writes_3_values_1 ^ writes_3_values_2));
  assign reads_0_values_0 = _zz_ram_0_port4;
  assign reads_0_values_1 = _zz_ram_1_port4;
  assign reads_0_values_2 = _zz_ram_2_port4;
  assign reads_0_values_3 = _zz_ram_3_port4;
  assign reads_0_xored = ((reads_0_values_0 ^ reads_0_values_1) ^ (reads_0_values_2 ^ reads_0_values_3));
  assign io_read_0_rsp = reads_0_xored;
  assign reads_1_values_0 = _zz_ram_0_port5;
  assign reads_1_values_1 = _zz_ram_1_port5;
  assign reads_1_values_2 = _zz_ram_2_port5;
  assign reads_1_values_3 = _zz_ram_3_port5;
  assign reads_1_xored = ((reads_1_values_0 ^ reads_1_values_1) ^ (reads_1_values_2 ^ reads_1_values_3));
  assign io_read_1_rsp = reads_1_xored;
  assign reads_2_values_0 = _zz_ram_0_port6;
  assign reads_2_values_1 = _zz_ram_1_port6;
  assign reads_2_values_2 = _zz_ram_2_port6;
  assign reads_2_values_3 = _zz_ram_3_port6;
  assign reads_2_xored = ((reads_2_values_0 ^ reads_2_values_1) ^ (reads_2_values_2 ^ reads_2_values_3));
  assign io_read_2_rsp = reads_2_xored;
  assign reads_3_values_0 = _zz_ram_0_port7;
  assign reads_3_values_1 = _zz_ram_1_port7;
  assign reads_3_values_2 = _zz_ram_2_port7;
  assign reads_3_values_3 = _zz_ram_3_port7;
  assign reads_3_xored = ((reads_3_values_0 ^ reads_3_values_1) ^ (reads_3_values_2 ^ reads_3_values_3));
  assign io_read_3_rsp = reads_3_xored;
  assign reads_4_values_0 = _zz_ram_0_port8;
  assign reads_4_values_1 = _zz_ram_1_port8;
  assign reads_4_values_2 = _zz_ram_2_port8;
  assign reads_4_values_3 = _zz_ram_3_port8;
  assign reads_4_xored = ((reads_4_values_0 ^ reads_4_values_1) ^ (reads_4_values_2 ^ reads_4_values_3));
  assign io_read_4_rsp = reads_4_xored;
  assign reads_5_values_0 = _zz_ram_0_port9;
  assign reads_5_values_1 = _zz_ram_1_port9;
  assign reads_5_values_2 = _zz_ram_2_port9;
  assign reads_5_values_3 = _zz_ram_3_port9;
  assign reads_5_xored = ((reads_5_values_0 ^ reads_5_values_1) ^ (reads_5_values_2 ^ reads_5_values_3));
  assign io_read_5_rsp = reads_5_xored;

endmodule
