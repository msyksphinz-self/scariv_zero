module msrh_ptw
  (
   // Page Table Walk I/O
   tlb_ptw_if.slave ptw_if
   );

endmodule // msrh_ptw
