package msrh_fpu_pkg;

import decoder_fpu_ctrl_pkg::*;

typedef struct packed {
  size_t size;
  op_t   op;
} pipe_ctrl_t;

endpackage // msrh_fpu_pkg
